/********************
* Filename:     bfm_arbiter.v
* Description:  Bus functional model to check the functionality of Arbiter which decides which of the Input port buffer gets the highest priority among the others. Arbitration is based on Round-Robin Scheduling policy with the last served as least priority. Priority direction Local, North, East, South, West
*
* $Revision: 26 $
* $Id: bfm_arbiter.v 26 2015-11-22 19:24:28Z ranga $
* $Date: 2015-11-22 21:24:28 +0200 (Sun, 22 Nov 2015) $
* $Author: ranga $
*********************/
`include "../DUTs/parameters.v"
`include "../DUTs/state_defines.v"

module bfm_arbiter(bfm_clk, bfm_command, bfm_grant);

  input bfm_clk;
  input [5:0] bfm_command;
  
  output reg bfm_grant;
  
  // Declaring the port variables for DUT
  wire        clk;
  
  reg         rst;
  reg [2:0]   Lflit_id, Nflit_id, Eflit_id, Wflit_id, Sflit_id;
  reg [11:0]  Llength, Nlength, Elength, Wlength, Slength;
  reg         Lreq, Nreq, Ereq, Wreq, Sreq;
  
  wire [5:0] nextstate;
  
  // Specifying timeout period
  parameter TIMEOUT = 5;
  integer loop;
  
  always @(negedge clk) begin
    if(!rst) begin
      {Lflit_id, Nflit_id, Eflit_id, Wflit_id, Sflit_id} = {`HEADER, `HEADER, `HEADER, `HEADER, `HEADER};
      Llength = TIMEOUT;
      Nlength = TIMEOUT;
      Elength = TIMEOUT;
      Wlength = TIMEOUT;
      Slength = TIMEOUT;
      for(loop = 0; loop < TIMEOUT-1; loop = loop + 1) begin
        @(negedge clk) begin
          {Lflit_id, Nflit_id, Eflit_id, Wflit_id, Sflit_id} = {`PAYLOAD, `PAYLOAD, `PAYLOAD, `PAYLOAD, `PAYLOAD};
        end
      end
      {Lflit_id, Nflit_id, Eflit_id, Wflit_id, Sflit_id} = {`TAIL, `TAIL, `TAIL, `TAIL, `TAIL};
    end
  end
  
  // Specifying the single pulse request parameter
  parameter NR = 3'b000,        // No request
            RS = 3'b001,        // Request to south
            RW = 3'b010,        // Request to west
            RE = 3'b011,        // Request to east
            RN = 3'b100,        // Request to north
            RL = 3'b101;        // Request to local
            
  // Specifying the continuous pulse(with access time) request parameter
  // Adding Extra bit for FSM Transition. To differentiate L-->N(00001), N-->L(10001). MSB stands for forward/backward
  parameter NRQ   = 6'b00000,           // No request
            RLN   = 6'b00001,           // Local to north
            RLE   = 6'b00010,           // Local to east
            RLW   = 6'b00011,           // Local to west
            RLS   = 6'b00100,           // Local to south
            RLL   = 6'b00101,           // Local to local
            RNE   = 6'b00110,           // North to east
            RNW   = 6'b00111,           // North to west
            RNS   = 6'b01000,           // North to south
            RNL   = 6'b10001,           // North to local
            RNN   = 6'b01001,           // North to north
            REW   = 6'b01010,           // East to west
            RES   = 6'b01011,           // East to south
            REL   = 6'b10010,           // East to local
            REN   = 6'b10110,           // East to north
            REE   = 6'b01100,           // East to east
            RWS   = 6'b01101,           // West to south
            RWL   = 6'b10011,           // West to local
            RWN   = 6'b10111,           // West to north
            RWE   = 6'b11010,           // West to east
            RWW   = 6'b01110,           // West to west
            RSL   = 6'b10100,           // South to local
            RSN   = 6'b11000,           // South to north
            RSE   = 6'b11011,           // South to east
            RSW   = 6'b11101,           // South to west
            RSS   = 6'b01111,           // South to south
            RNE_L = 6'b010000,          // North and East to Local 
            RNW_L = 6'b010001,          // North and West to Local 
            RNS_L = 6'b010010,          // North and South to Local 
            REW_L = 6'b010011,          // East and West to Local 
            RES_L = 6'b010100,          // East and South to Local 
            RWS_L = 6'b010101,          // West and South to Local 
            RLE_N = 6'b010110,          // Local and East to North
            RLW_N = 6'b010111,          // Local and West to North
            RLS_N = 6'b011000,          // Local and South to North
            REW_N = 6'b011001,          // East and West to North
            RES_N = 6'b011010,          // East and South to North
            RWS_N = 6'b011011,          // West and South to North
            RLN_E = 6'b011100,          // Local and North to East
            RLW_E = 6'b011101,          // Local and West to East
            RLS_E = 6'b011110,          // Local and South to East
            RNW_E = 6'b011111,          // North and West to East
            RNS_E = 6'b100000,          // North and South to East
            RWS_E = 6'b100001,          // West and South to East
            RLN_W = 6'b100010,          // Local and North to West
            RLE_W = 6'b100011,          // Local and East to West
            RLS_W = 6'b100100,          // Local and South to West
            RNE_W = 6'b100101,          // North and East to West
            RNS_W = 6'b100110,          // North and South to West
            RES_W = 6'b100111,          // East and South to West
            RLN_S = 6'b101000,          // Local and North to South
            RLE_S = 6'b101001,          // Local and East to South
            RLW_S = 6'b101010,          // Local and West to South
            RNE_S = 6'b101011,          // North and East to South
            RNW_S = 6'b101100,          // North and West to South
            REW_S = 6'b101101;          // East and West to South          
  
  // BFM commands Declaration
  parameter NOREQ1 = 6'd1,
            REQFL  = 6'd2,
            REQFN  = 6'd3,
            REQFE  = 6'd4,
            REQFW  = 6'd5,
            REQFS  = 6'd6,
            NOREQ2 = 6'd7,
            REQFLN = 6'd8,
            REQFLE = 6'd9,
            REQFLW = 6'd10,
            REQFLS = 6'd11,
            REQFLL = 6'd12,
            REQFNE = 6'd13,
            REQFNW = 6'd14,
            REQFNS = 6'd15,
            REQFNL = 6'd16,
            REQFNN = 6'd17,
            REQFEW = 6'd18,
            REQFES = 6'd19,
            REQFEL = 6'd20,
            REQFEN = 6'd21,
            REQFEE = 6'd22,
            REQFWS = 6'd23,
            REQFWL = 6'd24,
            REQFWN = 6'd25,
            REQFWE = 6'd26,
            REQFWW = 6'd27,
            REQFSL = 6'd28,
            REQFSN = 6'd29,
            REQFSE = 6'd30,
            REQFSW = 6'd31,
            REQFSS = 6'd32, 
            REQFNE_L = 6'd33, 
            REQFNW_L = 6'd34, 
            REQFNS_L = 6'd35, 
            REQFEW_L = 6'd36, 
            REQFES_L = 6'd37, 
            REQFWS_L = 6'd38,   
            REQFLE_N = 6'd39,
            REQFLW_N = 6'd40,
            REQFLS_N = 6'd41,
            REQFEW_N = 6'd42,
            REQFES_N = 6'd43,
            REQFWS_N = 6'd44,
            REQFLN_E = 6'd45,
            REQFLW_E = 6'd46,
            REQFLS_E = 6'd47,
            REQFNW_E = 6'd48,
            REQFNS_E = 6'd49,
            REQFWS_E = 6'd50,
            REQFLN_W = 6'd51,
            REQFLE_W = 6'd52,
            REQFLS_W = 6'd53,
            REQFNE_W = 6'd54,
            REQFNS_W = 6'd55,
            REQFES_W = 6'd56,
            REQFLN_S = 6'd57, 
            REQFLE_S = 6'd58, 
            REQFLW_S = 6'd59, 
            REQFNE_S = 6'd60, 
            REQFNW_S = 6'd61, 
            REQFEW_S = 6'd62;  

  assign clk = bfm_clk;
  
  // Instantiate ARBITER DUT              
  arbiter DUT (clk, rst,
                Lflit_id, Nflit_id, Eflit_id, Wflit_id, Sflit_id,
                Llength, Nlength, Elength, Wlength, Slength,
                Lreq, Nreq, Ereq, Wreq, Sreq,
                nextstate
              );
              
  // Task to generate reset
  task reset;
    begin
      rst                                                 = 1;
      {Lflit_id, Nflit_id, Eflit_id, Wflit_id, Sflit_id}  = 0;
      {Llength, Nlength, Elength, Wlength, Slength}       = 0;
      {Lreq, Nreq, Ereq, Wreq, Sreq}                      = 0;
      @(negedge clk);
        if(nextstate != `IDLE) begin
          $display("Reset is not working\n");
          $display("Error at time %0t", $time);
          $stop; 
        end
        $display("TIME:%0t Reset is working\n", $time);
        repeat(2)
          @(negedge clk);
        rst = 0;
    end
  endtask
  
  // Task to request buffer for first time -- single pulse
  task request1;
    input [2:0] data;
    begin
      @(negedge clk) begin
        if(data == 0) begin
          {Lreq, Nreq, Ereq, Wreq, Sreq} = 0;
        end
        else begin
          {Lreq, Nreq, Ereq, Wreq, Sreq} = (1 << (data-1)); // To assert the particular bit since data == 0 is used for IDLE
        end
      end
    end
  endtask
  
  // Task to request buffer for first time withoout last request -- continuous pulse requested by any buffer
  task request2;
    input Lr, Nr, Er, Wr, Sr;
    input [4:0] data;
    begin
      @(negedge clk) begin
        if(data == 0) begin
          {Lreq, Nreq, Ereq, Wreq, Sreq} = 0;
        end
        else begin
          {Lreq, Nreq, Ereq, Wreq, Sreq} = {Lr, Nr, Er, Wr, Sr};
        end
      end
      
      repeat(TIMEOUT+2) //Repeating the request for a particular buffer till timeout occurs followed by round robin priority request
        @(negedge clk);
    end
  endtask
  
  // Sampling and executing Commands
  always @(posedge clk) begin
    case(bfm_command)
      NOREQ1 :
        begin
          bfm_grant = 1'b0;
          request1(NR);
          bfm_grant = 1'b1;
        end
      REQFL :
        begin
          bfm_grant = 1'b0;
          request1(RL);
          request1(NR);
          bfm_grant = 1'b1;
        end
      REQFN :
        begin
          bfm_grant = 1'b0;
          request1(RN);
          request1(NR);
          bfm_grant = 1'b1;
        end
      REQFE :
        begin
          bfm_grant = 1'b0;
          request1(RE);
          request1(NR);
          bfm_grant = 1'b1;
        end
      REQFW :
        begin
          bfm_grant = 1'b0;
          request1(RW);
          request1(NR);
          bfm_grant = 1'b1;
        end
      REQFS :
        begin
          bfm_grant = 1'b0;
          request1(RS);
          request1(NR);
          bfm_grant = 1'b1;
        end
      NOREQ2 :
        begin
          bfm_grant = 1'b0;
          request2(0, 0, 0, 0, 0, NRQ);
          bfm_grant = 1'b1;
        end
      REQFLN :
        begin
          bfm_grant = 1'b0;
          request2(1, 1, 1, 1, 1, RLN);
          bfm_grant = 1'b1;
        end
      REQFLE :
        begin
          bfm_grant = 1'b0;
          request2(1, 0, 1, 1, 1, RLE);
          bfm_grant = 1'b1;
        end
      REQFLW :
        begin
          bfm_grant = 1'b0;
          request2(0, 0, 0, 1, 0, RLW);
          bfm_grant = 1'b1;
        end
      REQFLS :
        begin
          bfm_grant = 1'b0;
          request2(1, 0, 0, 0, 1, RLS);
          bfm_grant = 1'b1;
        end
      REQFLL :
        begin
          bfm_grant = 1'b0;
          request2(1, 0, 0, 0, 0, RLL);
          bfm_grant = 1'b1;
        end
      REQFNE :
        begin
          bfm_grant = 1'b0;
          request2(1, 1, 1, 1, 1, RNE);
          bfm_grant = 1'b1;
        end
      REQFNW :
        begin
          bfm_grant = 1'b0;
          request2(1, 1, 0, 1, 1, RNW);
          bfm_grant = 1'b1;
        end
      REQFNS :
        begin
          bfm_grant = 1'b0;
          request2(1, 1, 0, 0, 1, RNS);
          bfm_grant = 1'b1;
        end
      REQFNL :
        begin
          bfm_grant = 1'b0;
          request2(1, 0, 0, 0, 0, RNL);
          bfm_grant = 1'b1;
        end
      REQFNN :
        begin
          bfm_grant = 1'b0;
          request2(0, 1, 0, 0, 0, RNN);
          bfm_grant = 1'b1;
        end
      REQFEW :
        begin
          bfm_grant = 1'b0;
          request2(1, 1, 1, 1, 1, REW);
          bfm_grant = 1'b1;
        end
      REQFES :
        begin
          bfm_grant = 1'b0;
          request2(1, 1, 1, 0, 1, RES);
          bfm_grant = 1'b1;
        end
      REQFEL :
        begin
          bfm_grant = 1'b0;
          request2(1, 1, 1, 0, 0, REL);
          bfm_grant = 1'b1;
        end
      REQFEN :
        begin
          bfm_grant = 1'b0;
          request2(0, 1, 1, 0, 0, REN);
          bfm_grant = 1'b1;
        end
      REQFEE :
        begin
          bfm_grant = 1'b0;
          request2(0, 0, 1, 0, 0, REE);
          bfm_grant = 1'b1;
        end
      REQFWS :
        begin
          bfm_grant = 1'b0;
          request2(1, 1, 1, 1, 1, RWS);
          bfm_grant = 1'b1;
        end
      REQFWL :
        begin
          bfm_grant = 1'b0;
          request2(1, 1, 1, 1, 0, RWL);
          bfm_grant = 1'b1;
        end
      REQFWN :
        begin
          bfm_grant = 1'b0;
          request2(0, 1, 1, 1, 0, RWN);
          bfm_grant = 1'b1;
        end
      REQFWE :
        begin
          bfm_grant = 1'b0;
          request2(0, 0, 1, 1, 0, RWE);
          bfm_grant = 1'b1;
        end
      REQFWW :
        begin
          bfm_grant = 1'b0;
          request2(0, 0, 0, 1, 0, RWW);
          bfm_grant = 1'b1;
        end
      REQFSL :
        begin
          bfm_grant = 1'b0;
          request2(1, 0, 0, 0, 0, RSL);
          bfm_grant = 1'b1;
        end
      REQFSN :
        begin
          bfm_grant = 1'b0;
          request2(0, 1, 0, 0, 0, RSN);
          bfm_grant = 1'b1;
        end
      REQFSE :
        begin
          bfm_grant = 1'b0;
          request2(0, 0, 1, 0, 0, RSE);
          bfm_grant = 1'b1;
        end
      REQFSW :
        begin
          bfm_grant = 1'b0;
          request2(0, 0, 0, 1, 0, RSW);
          bfm_grant = 1'b1;
        end
      REQFSS :
        begin
          bfm_grant = 1'b0;
          request2(0, 0, 0, 0, 1, RSS);
          bfm_grant = 1'b1;
        end

      // Two requests to Local
      REQFNE_L :
        begin
          bfm_grant = 1'b0;
          request2(0, 1, 1, 0, 0, RNE_L);
          bfm_grant = 1'b1;
        end

      REQFNW_L :
        begin
          bfm_grant = 1'b0;
          request2(0, 1, 0, 1, 0, RNW_L);
          bfm_grant = 1'b1;
        end

      REQFNS_L :
        begin
          bfm_grant = 1'b0;
          request2(0, 1, 0, 0, 1, RNS_L);
          bfm_grant = 1'b1;
        end

      REQFEW_L :
        begin
          bfm_grant = 1'b0;
          request2(0, 0, 1, 1, 0, REW_L);
          bfm_grant = 1'b1;
        end

      REQFES_L :
        begin
          bfm_grant = 1'b0;
          request2(0, 0, 1, 0, 1, RES_L);
          bfm_grant = 1'b1;
        end

      REQFWS_L :
        begin
          bfm_grant = 1'b0;
          request2(0, 0, 0, 1, 1, RWS_L);
          bfm_grant = 1'b1;
        end
        
    endcase
  end

// Properties


property property_0;
@(negedge clk)
(rst) |->  nextstate[0];
endproperty

property property_1;
@(negedge clk)
 !Lreq && !Nreq && !Ereq && !Wreq && !Sreq |->  nextstate[0];
endproperty

property property_2;
@(negedge clk)
!rst && Lflit_id[2]  && Lreq && !Nreq && !Ereq && !Wreq && !Sreq |-> !nextstate[0];
endproperty

property property_3;
@(negedge clk)
 !rst && Lflit_id[2]  && Sreq |-> !nextstate[0];
endproperty

property property_4;
@(negedge clk)
 !rst && !Lflit_id[2]  && !Lflit_id[1] && !Nflit_id[2]  && !Eflit_id[2]  && !Wflit_id[2]  && !Sflit_id[2]  && Sreq |-> !nextstate[0];
endproperty

property property_5;
@(negedge clk)
 !rst && Lflit_id[0] && !Lreq && !Nreq && Ereq && !Sreq |-> !nextstate[0];
endproperty

property property_6;
@(negedge clk)
 !rst && Lflit_id[0] && !Lreq && !Nreq && !Ereq && Wreq && !Sreq |-> !nextstate[0];
endproperty

property property_7;
@(negedge clk)
 !rst && Lflit_id[0] && Nreq && !Sreq |-> !nextstate[0];
endproperty

property property_8;
@(negedge clk)
 !rst && !Lflit_id[0] && !Nflit_id[0] && !Eflit_id[0] && !Wflit_id[0] && !Sflit_id[0] && Lreq && Nreq && !Wreq && !Sreq |-> !nextstate[0];
endproperty

property property_9;
@(negedge clk)
 !rst && !Lflit_id[0] && !Nflit_id[0] && !Eflit_id[0] && !Wflit_id[0] && !Sflit_id[0] && !Lreq && Nreq && Ereq && !Wreq && !Sreq |-> !nextstate[0];
endproperty

property property_10;
@(negedge clk)
 !rst && !Lflit_id[0] && !Nflit_id[0] && !Eflit_id[0] && !Wflit_id[0] && !Sflit_id[0] && !Lreq && !Nreq && Ereq && Wreq && !Sreq |-> !nextstate[0];
endproperty

property property_11;
@(negedge clk)
 !rst && !Lflit_id[0] && !Nflit_id[0] && !Eflit_id[0] && !Wflit_id[0] && !Sflit_id[0] && Nreq && Wreq && !Sreq |-> !nextstate[0];
endproperty

property property_12;
@(negedge clk)
 !rst && !Lreq |-> !nextstate[1];
endproperty

property property_13;
@(negedge clk)
(rst) |-> !nextstate[1];
endproperty

property property_14;
@(negedge clk)
 Lflit_id[0] && !Lreq && Nreq && !Ereq |->  nextstate[2];
endproperty

property property_15;
@(negedge clk)
 Lflit_id[0] && Nreq && !Ereq && !Sreq |-> nextstate[2];
endproperty

property property_16;
@(negedge clk)
 !rst && Lflit_id[2]  && !Lflit_id[0] && !Nflit_id[0] && !Eflit_id[0] && !Wflit_id[0] && !Sflit_id[0] && Lreq && Nreq && !Wreq |-> !nextstate[2];
endproperty

property property_17;
@(negedge clk)
 !rst && Lflit_id[0] && Lreq && Nreq && !Wreq |-> !nextstate[2];
endproperty

property property_18;
@(negedge clk)
 !rst && !Nreq |-> !nextstate[2];
endproperty

property property_19;
@(negedge clk)
(rst) |-> !nextstate[2];
endproperty

property property_20;
@(negedge clk)
 Lflit_id[0] && !Nreq && Ereq && !Wreq |-> nextstate[3];
endproperty

property property_21;
@(negedge clk)
 !rst && Lflit_id[2]  && !Lreq && Nreq && Ereq && !Sreq |-> !nextstate[3];
endproperty

property property_22;
@(negedge clk)
 !rst && !Lflit_id[2]  && !Nflit_id[2]  && !Eflit_id[2]  && !Wflit_id[2]  && !Sflit_id[2]  && !Lreq && Nreq && Ereq && Wreq && !Sreq |-> !nextstate[3];
endproperty

property property_23;
@(negedge clk)
 !rst && !Ereq |-> !nextstate[3];
endproperty

property property_24;
@(negedge clk)
(rst) |-> !nextstate[3];
endproperty

property property_25;
@(negedge clk)
 !rst && !Wreq |-> !nextstate[4];
endproperty

property property_26;
@(negedge clk)
(rst) |-> !nextstate[4];
endproperty

property property_27;
@(negedge clk)
rst |-> nextstate[0];
endproperty

property property_28;
@(negedge clk)
 !rst && Lflit_id[2]  && !Lflit_id[0] && !Nflit_id[0] && !Eflit_id[0] && !Wflit_id[0] && !Sflit_id[0] && !Lreq && !Nreq && Ereq && !Sreq |-> ##1 !nextstate[0];
endproperty

property property_29;
@(negedge clk)
 !rst && Lflit_id[2]  && !Lreq && !Nreq && !Ereq && Wreq && !Sreq |-> ##1  !nextstate[0];
endproperty

property property_30;
@(negedge clk)
 !rst && Lflit_id[2]  && Sreq |-> ##1 !nextstate[0];
endproperty

property property_31;
@(negedge clk)
 !rst && !Lflit_id[2]  && !Nflit_id[2]  && !Eflit_id[2]  && !Wflit_id[2]  && !Sflit_id[2]  && Lreq && !Nreq && !Ereq && !Wreq && Sreq |-> ##1 !nextstate[0];
endproperty

property property_32;
@(negedge clk)
 !rst && !Lflit_id[2]  && !Nflit_id[2]  && !Eflit_id[2]  && !Wflit_id[2]  && !Sflit_id[2]  && Nreq && !Ereq && !Wreq && Sreq |-> ##1 !nextstate[0];
endproperty

property property_33;
@(negedge clk)
 !rst && !Lflit_id[2]  && !Nflit_id[2]  && !Eflit_id[2]  && !Wflit_id[2]  && !Sflit_id[2]  && Ereq && Sreq |-> ##1 !nextstate[0];
endproperty

property property_34;
@(negedge clk)
 !rst && !Lflit_id[2]  && !Nflit_id[2]  && !Eflit_id[2]  && !Wflit_id[2]  && !Sflit_id[2]  && !Ereq && Wreq && Sreq |-> ##1 !nextstate[0];
endproperty

property property_35;
@(negedge clk)
 !rst && Lflit_id[0] && Lreq && !Nreq && !Ereq && !Wreq && !Sreq |-> ##1 !nextstate[0];
endproperty

property property_36;
@(negedge clk)
 !rst && Lflit_id[0] && !Lreq && !Nreq && Ereq && !Sreq |-> ##1 !nextstate[0];
endproperty

property property_37;
@(negedge clk)
 !rst && Lflit_id[0] && Nreq && Ereq && !Wreq && !Sreq |-> ##1 !nextstate[0];
endproperty

property property_38;
@(negedge clk)
 !rst && !Lflit_id[0] && !Nflit_id[0] && !Eflit_id[0] && !Wflit_id[0] && !Sflit_id[0] && !Lreq && Nreq && Ereq && !Wreq && !Sreq |-> ##1 !nextstate[0];
endproperty

property property_39;
@(negedge clk)
 !rst && Nreq && Wreq && !Sreq |-> ##1 !nextstate[0];
endproperty

property property_40;
@(negedge clk)
 !rst && Lflit_id[2]  && !Lflit_id[0] && !Nflit_id[0] && !Eflit_id[0] && !Wflit_id[0] && !Sflit_id[0] && Lreq && Nreq && !Wreq && !Sreq |-> ##1 !nextstate[1];
endproperty

property property_41;
@(negedge clk)
 !rst && Lflit_id[2]  && !Lflit_id[0] && !Nflit_id[0] && !Eflit_id[0] && !Wflit_id[0] && !Sflit_id[0] && !Lreq && Nreq && !Wreq && !Sreq |-> ##1 !nextstate[1];
endproperty

property property_42;
@(negedge clk)
 !rst && !Lflit_id[2]  && !Lflit_id[1] && !Nflit_id[2]  && !Eflit_id[2]  && !Wflit_id[2]  && !Sflit_id[2]  && Lreq && !Ereq && Sreq |-> ##1 !nextstate[1];
endproperty

property property_43;
@(negedge clk)
 !rst && !Lflit_id[2]  && !Nflit_id[2]  && !Eflit_id[2]  && !Wflit_id[2]  && !Sflit_id[2]  && Lreq && !Nreq && Ereq && Sreq |-> ##1 !nextstate[1];
endproperty

property property_44;
@(negedge clk)
 !rst && Lflit_id[0] && !Lreq && !Sreq |-> ##1 !nextstate[1];
endproperty

property property_45;
@(negedge clk)
 !rst && !Lflit_id[0] && !Nflit_id[0] && !Eflit_id[0] && !Wflit_id[0] && !Sflit_id[0] && !Lreq && !Nreq && Ereq && !Wreq && !Sreq |-> ##1 !nextstate[1];
endproperty

property property_46;
@(negedge clk)
 !rst && !Lflit_id[0] && !Nflit_id[0] && !Eflit_id[0] && !Wflit_id[0] && !Sflit_id[0] && !Lreq && Wreq && !Sreq |-> ##1 !nextstate[1];
endproperty

property property_47;
@(negedge clk)
 !rst && !Lreq && Sreq |-> ##1 !nextstate[1];
endproperty

property property_48;
@(negedge clk)
(rst) |-> ##1 !nextstate[1];
endproperty

property property_49;
@(negedge clk)
 !rst && Lflit_id[2]  && !Lflit_id[0] && !Nflit_id[0] && !Eflit_id[0] && !Wflit_id[0] && !Sflit_id[0] && Lreq && Nreq && !Wreq |-> ##1 !nextstate[2];
endproperty

property property_50;
@(negedge clk)
 !rst && Lflit_id[2]  && !Nreq |-> ##1 !nextstate[2];
endproperty

property property_51;
@(negedge clk)
 !rst && !Lflit_id[2]  && !Lflit_id[1] && !Nflit_id[2]  && !Eflit_id[2]  && !Wflit_id[2]  && !Sflit_id[2]  && !Nreq && !Ereq && !Sreq |-> ##1 !nextstate[2];
endproperty

property property_52;
@(negedge clk)
 !rst && !Lflit_id[2]  && !Nflit_id[2]  && !Eflit_id[2]  && !Wflit_id[2]  && !Sflit_id[2]  && !Nreq && Ereq && !Sreq |-> ##1 !nextstate[2];
endproperty

property property_53;
@(negedge clk)
 !rst && !Lflit_id[2]  && !Nflit_id[2]  && !Eflit_id[2]  && !Wflit_id[2]  && !Sflit_id[2]  && !Nreq && Sreq |-> ##1 !nextstate[2];
endproperty

property property_54;
@(negedge clk)
 !rst && Lflit_id[0] && Lreq && Nreq && Ereq && Wreq && !Sreq |-> ##1 !nextstate[2];
endproperty

property property_55;
@(negedge clk)
 !rst && Lflit_id[0] && Lreq && Nreq && !Wreq |-> ##1 !nextstate[2];
endproperty

property property_56;
@(negedge clk)
(rst) |-> ##1 !nextstate[2];
endproperty

property property_57;
@(negedge clk)
 Lflit_id[0] && !Nreq && Ereq && !Wreq |-> ##1 nextstate[3];
endproperty

property property_58;
@(negedge clk)
 !rst && Lflit_id[2]  && !Lreq && Nreq && Ereq && !Sreq |-> ##1 !nextstate[3];
endproperty

property property_59;
@(negedge clk)
 !rst && Lflit_id[2]  && !Ereq |-> ##1 !nextstate[3];
endproperty

property property_60;
@(negedge clk)
 !rst && !Lflit_id[2]  && !Lflit_id[1]&& !Nflit_id[2]  && !Eflit_id[2]  && !Wflit_id[2]  && !Sflit_id[2]  && Lreq && !Ereq && !Wreq |-> ##1 !nextstate[3];
endproperty

property property_61;
@(negedge clk)
 !rst && !Lflit_id[2]  && !Lflit_id[1]&& !Nflit_id[2]  && !Eflit_id[2]  && !Wflit_id[2]  && !Sflit_id[2]  && !Lreq && Nreq && Ereq && !Sreq |-> ##1 !nextstate[3];
endproperty

property property_62;
@(negedge clk)
 !rst && !Lflit_id[2]  && !Lflit_id[1]&& !Nflit_id[1] && !Eflit_id[1] && !Wflit_id[1] && !Sflit_id[2]  && Lreq && Nreq && Ereq && !Sreq |-> ##1 !nextstate[3];
endproperty

property property_63;
@(negedge clk)
 !rst && !Lflit_id[2]  && !Nflit_id[2]  && !Eflit_id[2]  && !Wflit_id[2]  && !Sflit_id[2]  && !Lreq && Nreq && !Ereq && !Wreq && !Sreq |-> ##1 !nextstate[3];
endproperty

property property_64;
@(negedge clk)
 !rst && !Lflit_id[2]  && !Nflit_id[2]  && !Eflit_id[2]  && !Wflit_id[2]  && !Sflit_id[2]  && !Lreq && !Ereq && !Wreq && Sreq |-> ##1 !nextstate[3];
endproperty

property property_65;
@(negedge clk)
 !rst && !Lflit_id[2]  && !Nflit_id[2]  && !Eflit_id[2]  && !Wflit_id[2]  && !Sflit_id[2]  && !Ereq && Wreq |-> ##1 !nextstate[3];
endproperty

property property_66;
@(negedge clk)
 !rst && !Lflit_id[1] && !Nflit_id[1] && !Eflit_id[1] && !Wflit_id[1] && !Sflit_id[2]  && Lreq && Nreq && Ereq && !Wreq && Sreq |-> ##1 !nextstate[3];
endproperty

property property_67;
@(negedge clk)
(rst) |-> ##1 !nextstate[3];
endproperty

property property_68;
@(negedge clk)
 Lflit_id[2]  && !Ereq && Wreq |-> ##1 nextstate[4];
endproperty

property property_69;
@(negedge clk)
 !rst && Lflit_id[2]  && !Wreq |-> ##1 !nextstate[4];
endproperty

property property_70;
@(negedge clk)
 !rst && !Lflit_id[2]  && !Lflit_id[1] && !Nflit_id[2]  && !Eflit_id[2]  && !Wflit_id[2]  && !Sflit_id[2]  && !Wreq |-> ##1 !nextstate[4];
endproperty

property property_71;
@(negedge clk)
 !rst && !Lflit_id[0] && !Nflit_id[0] && !Eflit_id[0] && !Wflit_id[0] && !Sflit_id[0] && Lreq && Ereq && Wreq && !Sreq |-> ##1 !nextstate[4];
endproperty

property property_72;
@(negedge clk)
(rst) |-> ##1 !nextstate[4];
endproperty

property property_76;
@(negedge clk)
 !rst && Lflit_id[2]  && !Lreq && !Nreq && Ereq && !Sreq ##1 !rst && !Lreq && !Nreq && Ereq && !Sreq |-> ##1 !nextstate[0];
endproperty

property property_77;
@(negedge clk)
 !rst && Lflit_id[2] && Nreq && !Sreq ##1 !rst && Nreq && !Sreq |-> !nextstate[0];
endproperty

property property_79;
@(negedge clk)
 !rst && Lreq  ##1 !rst && !Lreq && !Nreq && Ereq && !Sreq |-> ##1 !nextstate[0];
endproperty

property property_80;
@(negedge clk)
 !rst && Lreq  ##1 !rst && !Lreq && !Nreq && !Ereq && Wreq && !Sreq |-> ##1 !nextstate[0];
endproperty

property property_82;
@(negedge clk)
 !rst && !Lreq && !Nreq && !Ereq && Sreq ##1 !rst && !Lreq && !Nreq && !Ereq && Wreq && !Sreq |-> ##1 !nextstate[0];
endproperty

property property_83;
@(negedge clk)
 !rst && Nreq && !Wreq && !Sreq  ##1 !rst && Lreq && !Nreq && !Ereq && !Wreq && !Sreq |-> ##1 !nextstate[0];
endproperty

property property_84;
@(negedge clk)
 !rst && Wreq  ##1 !rst && Lreq && !Nreq && !Ereq && !Wreq && !Sreq |-> ##1 !nextstate[0];
endproperty

property property_86;
@(negedge clk)
 !rst && Sreq ##1 !rst && Nreq && !Sreq |-> ##1 !nextstate[0];
endproperty

property property_92;
@(negedge clk)
rst ##1 !rst |-> ##1 !nextstate[1];
endproperty

property property_93;
@(negedge clk)
Lreq ##1  !Lreq && Nreq |-> ##1  nextstate[2];
endproperty

property property_96;
@(negedge clk)
 !rst && !Nreq ##1 !rst && Lreq && Nreq |-> ##1 !nextstate[2];
endproperty

property property_98;
@(negedge clk)
1 ##1 rst |-> ##1 !nextstate[2];
endproperty

property property_99;
@(negedge clk)
rst ##1 !rst |-> ##1 !nextstate[2];
endproperty

property property_100;
@(negedge clk)
 !Lreq && Ereq ##1  Lreq && Ereq |-> ##1  nextstate[3];
endproperty
property property_102;
@(negedge clk)
Nreq ##1 !Nreq && Ereq |-> ##1  nextstate[3];
endproperty

property property_103;
@(negedge clk)
 !rst && !Lreq && Nreq && Ereq && !Sreq ##1 !rst && Lflit_id[2]  && !Lreq && Nreq && Ereq && !Sreq |-> ##1 !nextstate[3];
endproperty

property property_105;
@(negedge clk)
 !rst && Lreq && !Nreq && Ereq  ##1 !rst && Lreq && Nreq && Ereq |-> ##1 !nextstate[3];
endproperty

property property_106;
@(negedge clk)
 !rst && !Ereq ##1 !rst && Nreq && Ereq |-> ##1 !nextstate[3];
endproperty

property property_108;
@(negedge clk)
1 ##1 rst |-> ##1 !nextstate[3];
endproperty

property property_109;
@(negedge clk)
rst ##1 !rst |-> ##1 !nextstate[3];
endproperty

property property_112;
@(negedge clk)
Ereq ##1  !Ereq && Wreq |-> ##1  nextstate[4];
endproperty

property property_114;
@(negedge clk)
 !rst && Lflit_id[2]  && !Ereq && !Wreq ##1 !rst && !Ereq && Wreq |-> ##1 !nextstate[4];
endproperty

property property_115;
@(negedge clk)
 !rst && !Wreq ##1 !rst && Ereq && Wreq |-> ##1 !nextstate[4];
endproperty

property property_117;
@(negedge clk)
1 ##1 rst |-> ##1 !nextstate[4];
endproperty

property property_118;
@(negedge clk)
rst ##1 !rst |-> ##1 !nextstate[4];
endproperty

property property_121;
@(negedge clk)
 !Lflit_id[1] && Sreq ##1 !Sreq |-> ##1  nextstate[0];
endproperty

property property_122;
@(negedge clk)
 Lreq && Nreq && !Wreq && !Sreq ##1 !Nreq |-> ##1  nextstate[0];
endproperty

property property_123;
@(negedge clk)
 !Lreq && !Nreq ##1  Lreq && !Nreq |-> ##1  nextstate[0];
endproperty

property property_124;
@(negedge clk)
 !Lreq && !Ereq ##1  Lreq && !Nreq |-> ##1  nextstate[0];
endproperty

property property_125;
@(negedge clk)
 !Lreq && !Ereq && !Wreq ##1  !Lreq && Ereq |-> ##1  nextstate[0];
endproperty

property property_126;
@(negedge clk)
 !Lreq && !Ereq && !Wreq ##1 !Nreq && Ereq |-> ##1  nextstate[0];
endproperty

property property_127;
@(negedge clk)
 !Nreq && !Ereq && !Wreq ##1  !Lreq && Ereq |-> ##1  nextstate[0];
endproperty

property property_128;
@(negedge clk)
 !Ereq && !Wreq && !Sreq ##1  !Lreq && Ereq |-> ##1  nextstate[0];
endproperty

property property_129;
@(negedge clk)
 !Wreq && !Sreq ##1  !Lreq && Wreq |-> ##1  nextstate[0];
endproperty

property property_130;
@(negedge clk)
 !rst && !Lreq && !Nreq && Wreq && !Sreq ##1 !rst && Lflit_id[2]  && !Lreq && !Nreq && Wreq && !Sreq |-> ##1 !nextstate[0];
endproperty

property property_131;
@(negedge clk)
 !rst && Sreq ##1 !rst && Lflit_id[2] |-> ##1 !nextstate[0];
endproperty

property property_132;
@(negedge clk)
 !rst && Lflit_id[1] && Sreq ##1 !rst && !Lflit_id[2]  && !Nflit_id[2]  && !Eflit_id[2]  && !Wflit_id[2]  && !Sflit_id[2] |-> ##1 !nextstate[0];
endproperty

property property_133;
@(negedge clk)
 !rst && Lflit_id[0] && !Wreq && !Sreq ##1 !rst && Nreq && !Wreq && !Sreq |-> ##1 !nextstate[0];
endproperty

property property_134;
@(negedge clk)
 !rst && Lreq && !Nreq && !Ereq && !Wreq && !Sreq ##1 !rst && Lreq && !Nreq && Ereq |-> ##1 !nextstate[0];
endproperty

property property_135;
@(negedge clk)
 !rst && Lreq && !Nreq && !Ereq && !Wreq && !Sreq ##1 !rst && !Lreq && !Nreq |-> ##1 !nextstate[0];
endproperty

property property_136;
@(negedge clk)
 !rst && Lreq && Wreq && !Sreq ##1 !rst && !Lreq && Wreq && !Sreq |-> ##1 !nextstate[0];
endproperty

property property_137;
@(negedge clk)
 !rst && !Lreq && Nreq && Wreq && !Sreq ##1 !rst && !Lreq && Wreq && !Sreq |-> ##1 !nextstate[0];
endproperty

property property_138;
@(negedge clk)
 !rst && !Lreq && !Nreq && Wreq && !Sreq ##1 !rst && !Lreq && Nreq && Wreq && !Sreq |-> ##1 !nextstate[0];
endproperty

property property_139;
@(negedge clk)
 !rst && !Lreq && Nreq && !Wreq && !Sreq ##1 !rst && !Nreq |-> ##1 !nextstate[0];
endproperty

property property_140;
@(negedge clk)  
!rst && Wreq && !Sreq  ##1 !rst && Lreq && Wreq && !Sreq |-> ##1 !nextstate[0];
endproperty

property property_141;
@(negedge clk)
 !rst && !Wreq && !Sreq  ##1 !rst && Nreq && Wreq |-> ##1 !nextstate[0];
endproperty

property property_142;
@(negedge clk)
 !rst && Wreq && !Sreq  ##1 !rst && !Wreq && !Sreq |-> ##1 !nextstate[0];
endproperty

property property_143;
@(negedge clk)
 !rst && Wreq && !Sreq  ##1 !rst && Sreq |-> ##1 !nextstate[0];
endproperty

property property_144;
@(negedge clk)
!Lreq ##1 Ereq && Sreq |-> ##1  nextstate[1];
endproperty

property property_145;
@(negedge clk)
Sreq ##1  Lreq && !Sreq |-> ##1  nextstate[1];
endproperty

property property_146;
@(negedge clk)
 !rst && Lflit_id[2]  && !Lreq && !Sreq ##1 !rst && !Lreq && !Sreq |-> ##1 !nextstate[1];
endproperty

property property_147;
@(negedge clk)
 !rst && Ereq ##1 !rst && !Lflit_id[2]  && !Nflit_id[2]  && !Eflit_id[2]  && !Wflit_id[2]  && !Sflit_id[2]  && Lreq && !Ereq && Sreq |-> ##1 !nextstate[1];
endproperty

property property_148;
@(negedge clk)
 !rst && Lreq ##1 !rst && !Lreq |-> ##1 !nextstate[1];
endproperty

property property_149;
@(negedge clk)
 !rst && !Lreq && Sreq ##1 !rst && !Lreq && !Sreq |-> ##1 !nextstate[1];
endproperty

property property_150;
@(negedge clk)
 !rst && !Lreq ##1 !rst && !Lreq && Sreq |-> ##1 !nextstate[1];
endproperty

property property_152;
@(negedge clk)
rst ##1 !rst |-> ##1 !nextstate[1];
endproperty

property property_153;
@(negedge clk)
 Lreq ##1  !Lreq && Nreq |-> ##1  nextstate[2];
endproperty

property property_154;
@(negedge clk)
 !Lreq && Nreq ##1  Lreq && Wreq |-> ##1  nextstate[2];
endproperty

property property_155;
@(negedge clk)
 !rst && Lflit_id[2]  && Lreq && Nreq && !Wreq ##1 !rst && Lreq && Nreq && !Wreq |-> ##1 !nextstate[2];
endproperty

property property_156;
@(negedge clk)
 !rst && Lflit_id[2]  && !Nreq ##1 !rst && !Nreq |-> ##1 !nextstate[2];
endproperty

property property_157;
@(negedge clk)
 !rst && !Lflit_id[2]  && !Lreq && !Nreq && !Sreq ##1 !rst && !Lreq && Nreq && !Sreq |-> ##1 !nextstate[2];
endproperty

property property_158;
@(negedge clk)
 !rst && !Lreq && Nreq ##1 !rst && Lreq && Nreq && !Wreq |-> ##1 !nextstate[2];
endproperty

property property_159;
@(negedge clk)
 !rst && !Nreq ##1 !rst && Lreq && Nreq |-> ##1 !nextstate[2];
endproperty

property property_160;
@(negedge clk)
 !rst && Nreq ##1 !rst && !Nreq |-> ##1 !nextstate[2];
endproperty

property property_162;
@(negedge clk)
rst ##1 !rst |-> ##1 !nextstate[2];
endproperty

property property_163;
@(negedge clk)
Lreq && !Nreq && !Wreq ##1 Ereq |-> ##1  nextstate[3];
endproperty

property property_164;
@(negedge clk)
Lreq && !Nreq && !Sreq ##1 Ereq |-> ##1  nextstate[3];
endproperty

property property_165;
@(negedge clk)
 Lreq && !Wreq ##1  !Nreq && Ereq |-> ##1  nextstate[3];
endproperty

property property_166;
@(negedge clk)
 Lreq && !Sreq ##1  !Nreq && Ereq |-> ##1  nextstate[3];
endproperty

property property_167;
@(negedge clk)
 !Lreq && Ereq ##1  Lreq && Ereq |-> ##1  nextstate[3];
endproperty

property property_168;
@(negedge clk)
Nreq ##1  !Nreq && Ereq |-> ##1  nextstate[3];
endproperty

property property_169;
@(negedge clk)
Wreq ##1  !Nreq && Ereq && !Wreq |-> ##1  nextstate[3];
endproperty

property property_170;
@(negedge clk)
 !rst && Lflit_id[2]  && !Lreq && Nreq && Ereq && !Sreq ##1 !rst && !Lreq && Nreq && Ereq && !Sreq |-> ##1 !nextstate[3];
endproperty

property property_171;
@(negedge clk)
 !rst && !Ereq ##1 !rst && Lflit_id[2]  && !Ereq |-> ##1 !nextstate[3];
endproperty

property property_172;
@(negedge clk)
 !rst && !Ereq && Wreq ##1 !rst && !Lflit_id[2]  && !Nflit_id[2]  && !Eflit_id[2]  && !Wflit_id[2]  && !Sflit_id[2]  && !Ereq |-> ##1 !nextstate[3];
endproperty

property property_173;
@(negedge clk)
 !rst && !Ereq && !Wreq ##1 !rst && !Lflit_id[2]  && !Nflit_id[2]  && !Eflit_id[2]  && !Wflit_id[2]  && !Sflit_id[2]  && !Ereq && Wreq |-> ##1 !nextstate[3];
endproperty

property property_174;
@(negedge clk)
 !rst && Lreq && !Nreq && Ereq ##1 !rst && Lreq && Nreq && Ereq |-> ##1 !nextstate[3];
endproperty

property property_175;
@(negedge clk)
 !rst && !Lreq && !Nreq && Ereq && !Sreq ##1 !rst && !Lreq && Nreq && Ereq && !Sreq |-> ##1 !nextstate[3];
endproperty

property property_176;
@(negedge clk)
 !rst && !Lreq && !Nreq && !Ereq && !Wreq && !Sreq ##1 !rst && !Nreq && Ereq |-> ##1 !nextstate[3];
endproperty

property property_177;
@(negedge clk)
 !rst && !Nreq && !Ereq && Wreq ##1 !rst && !Nreq && Ereq |-> ##1 !nextstate[3];
endproperty

property property_178;
@(negedge clk)
 !rst && !Ereq ##1 !rst && Nreq && Ereq |-> ##1 !nextstate[3];
endproperty

property property_179;
@(negedge clk)
 !rst && Ereq ##1 !rst && !Ereq |-> ##1 !nextstate[3];
endproperty

property property_180;
@(negedge clk)
1 ##1 rst |-> ##1 !nextstate[3];
endproperty

property property_181;
@(negedge clk)
rst ##1 !rst |-> ##1 !nextstate[3];
endproperty

property property_182;
@(negedge clk)
!Ereq ##1  Lflit_id[2]  && Wreq |-> ##1  nextstate[4];
endproperty

property property_183;
@(negedge clk)
1 ##1  Lflit_id[2]  && !Ereq && Wreq |-> ##1  nextstate[4];
endproperty

property property_184;
@(negedge clk)
 !Ereq && Wreq ##1  !Lflit_id[1] && Ereq |-> ##1  nextstate[4];
endproperty

property property_185;
@(negedge clk)
Ereq ##1  !Ereq && Wreq |-> ##1  nextstate[4];
endproperty

property property_186;
@(negedge clk)
 !rst && Lflit_id[2]  && !Wreq ##1 !rst && !Wreq |-> ##1 !nextstate[4];
endproperty

property property_187;
@(negedge clk)
 !rst && !Wreq ##1 !rst && Ereq && Wreq |-> ##1 !nextstate[4];
endproperty

property property_188;
@(negedge clk)
 !rst && Wreq ##1 !rst && !Wreq |-> ##1 !nextstate[4];
endproperty

property property_190;
@(negedge clk)
rst ##1 !rst |-> ##1 !nextstate[4];
endproperty


property property_n0; 
@(negedge clk)
!Sreq && !Wreq  &&   !Ereq  &&   !Nreq  &&   !Lreq |->  (nextstate[0]);
endproperty

property property_n1; 
@(negedge clk)
 rst |-> (nextstate[0]);
endproperty

property property_n2; 
@(negedge clk)
Sreq && Wreq  &&   !Nflit_id[2]  &&   !Sflit_id[0]  &&   Sflit_id[1] &&   !Sflit_id[2]  &&   !Wflit_id[0]  &&   Wflit_id[1] &&   !Wflit_id[2]  &&   !Eflit_id[0]  &&   Eflit_id[1] &&   !Eflit_id[2]  &&   !Nflit_id[0]  &&   Nflit_id[1] &&   !Lflit_id[0]  &&   Lflit_id[1] &&   !Lflit_id[2]  &&   !rst |->  (!nextstate[0]);
endproperty

property property_n3; 
@(negedge clk)
Sreq && !Wreq  &&   Ereq  &&   !Nflit_id[2]  &&   !Sflit_id[0]  &&   Sflit_id[1] &&   !Sflit_id[2]  &&   !Wflit_id[0]  &&   Wflit_id[1] &&   !Wflit_id[2]  &&   !Eflit_id[0]  &&   Eflit_id[1] &&   !Eflit_id[2]  &&   !Nflit_id[0]  &&   Nflit_id[1] &&   !Lflit_id[0]  &&   Lflit_id[1] &&   !Lflit_id[2]  &&   !rst |->  (!nextstate[0]);
endproperty

property property_n4; 
@(negedge clk)
Sreq && !Wreq  &&   !Ereq  &&   Nreq  &&   !Nflit_id[2]  &&   !Sflit_id[0]  &&   Sflit_id[1] &&   !Sflit_id[2]  &&   !Wflit_id[0]  &&   Wflit_id[1] &&   !Wflit_id[2]  &&   !Eflit_id[0]  &&   Eflit_id[1] &&   !Eflit_id[2]  &&   !Nflit_id[0]  &&   Nflit_id[1] &&   !Lflit_id[0]  &&   Lflit_id[1] &&   !Lflit_id[2]  &&   !rst |->  (!nextstate[0]);
endproperty

property property_n5; 
@(negedge clk)
Sreq && !Wreq  &&   !Ereq  &&   !Nreq  &&   Lreq  &&   !Nflit_id[2]  &&   !Sflit_id[0]  &&   Sflit_id[1] &&   !Sflit_id[2]  &&   !Wflit_id[0]  &&   Wflit_id[1] &&   !Wflit_id[2]  &&   !Eflit_id[0]  &&   Eflit_id[1] &&   !Eflit_id[2]  &&   !Nflit_id[0]  &&   Nflit_id[1] &&   !Lflit_id[0]  &&   Lflit_id[1] &&   !Lflit_id[2]  &&   !rst |->  (!nextstate[0]);
endproperty

property property_n6; 
@(negedge clk)
Sreq && !Nflit_id[2]  &&   !Sflit_id[2]  &&   !Wflit_id[2]  &&   !Eflit_id[2]  &&   !Lflit_id[1] &&   !Lflit_id[2]  &&   !rst |->  (!nextstate[0]);
endproperty

property property_n7; 
@(negedge clk)
Sreq && Lflit_id[2]  &&   !rst |->  (!nextstate[0]);
endproperty

property property_n8; 
@(negedge clk)
!Sreq && Wreq  &&   Ereq  &&   !Nreq  &&   !Lreq  &&   !Sflit_id[0]  &&   !Wflit_id[0]  &&   !Eflit_id[0]  &&   !Nflit_id[0]  &&   !Lflit_id[0]  &&   !rst |->  (!nextstate[0]);
endproperty

property property_n9; 
@(negedge clk)
!Sreq && Wreq  &&   !Ereq  &&   !Nreq  &&   !Lreq  &&   Lflit_id[0]  &&   !rst |->  (!nextstate[0]);
endproperty

property property_n10; 
@(negedge clk)
!Sreq && Wreq  &&   Nreq  &&   !Sflit_id[0]  &&   !Wflit_id[0]  &&   !Eflit_id[0]  &&   !Nflit_id[0]  &&   !Lflit_id[0]  &&   !rst |->  (!nextstate[0]);
endproperty

property property_n11; 
@(negedge clk)
!Sreq && !Wreq  &&   Ereq  &&   Nreq  &&   !Lreq  &&   !Sflit_id[0]  &&   !Wflit_id[0]  &&   !Eflit_id[0]  &&   !Nflit_id[0]  &&   !Lflit_id[0]  &&   !rst |->  (!nextstate[0]);
endproperty

property property_n12; 
@(negedge clk)
!Sreq && !Wreq  &&   Ereq  &&   !Nreq  &&   !Lreq  &&   !Sflit_id[0]  &&   !Wflit_id[0]  &&   !Eflit_id[0]  &&   !Nflit_id[0]  &&   !Lflit_id[0]  &&   !Lflit_id[2]  &&   !rst |->  (!nextstate[0]);
endproperty

property property_n13; 
@(negedge clk)
!Sreq && !Wreq  &&   !Ereq  &&   !Nreq  &&   Lreq  &&   Lflit_id[2]  &&   !rst |->  (!nextstate[0]);
endproperty

property property_n14; 
@(negedge clk)
!Sreq && !Wreq  &&   Nreq  &&   Lreq  &&   !Sflit_id[0]  &&   !Wflit_id[0]  &&   !Eflit_id[0]  &&   !Nflit_id[0]  &&   !Lflit_id[0]  &&   !rst |->  (!nextstate[0]);
endproperty

property property_n15; 
@(negedge clk)
!Sreq && Ereq  &&   !Nreq  &&   !Lreq  &&   Lflit_id[0]  &&   !rst |->  (!nextstate[0]);
endproperty

property property_n16; 
@(negedge clk)
!Sreq && Nreq  &&   Lflit_id[0]  &&   !rst |->  (!nextstate[0]);
endproperty

property property_n17; 
@(negedge clk)
!Sreq && Wreq  &&   Lreq  &&   Nflit_id[2] |->  (nextstate[1]);
endproperty

property property_n18; 
@(negedge clk)
!Sreq && Wreq  &&   Lreq  &&   Sflit_id[2] |->  (nextstate[1]);
endproperty

property property_n19; 
@(negedge clk)
!Sreq && Wreq  &&   Lreq  &&   Wflit_id[2] |->  (nextstate[1]);
endproperty

property property_n20; 
@(negedge clk)
!Sreq && Wreq  &&   Lreq  &&   Eflit_id[2] |->  (nextstate[1]);
endproperty

property property_n21; 
@(negedge clk)
!Sreq && Wreq  &&   Lreq  &&   Lflit_id[2] |->  (nextstate[1]);
endproperty

property property_n22; 
@(negedge clk)
!Sreq && !Nreq  &&   Lreq  &&   Nflit_id[2] |->  (nextstate[1]);
endproperty

property property_n23; 
@(negedge clk)
!Sreq && !Nreq  &&   Lreq  &&   Sflit_id[2] |->  (nextstate[1]);
endproperty

property property_n24; 
@(negedge clk)
!Sreq && !Nreq  &&   Lreq  &&   Wflit_id[2] |->  (nextstate[1]);
endproperty

property property_n25; 
@(negedge clk)
!Sreq && !Nreq  &&   Lreq  &&   Eflit_id[2] |->  (nextstate[1]);
endproperty

property property_n26; 
@(negedge clk)
!Sreq && !Nreq  &&   Lreq  &&   Lflit_id[2] |->  (nextstate[1]);
endproperty

property property_n27; 
@(negedge clk)
!Wreq && !Nreq  &&   Lreq  &&   Nflit_id[2] |->  (nextstate[1]);
endproperty

property property_n28; 
@(negedge clk)
!Wreq && !Nreq  &&   Lreq  &&   Sflit_id[2] |->  (nextstate[1]);
endproperty

property property_n29; 
@(negedge clk)
!Wreq && !Nreq  &&   Lreq  &&   Wflit_id[2] |->  (nextstate[1]);
endproperty

property property_n30; 
@(negedge clk)
!Wreq && !Nreq  &&   Lreq  &&   Eflit_id[2] |->  (nextstate[1]);
endproperty

property property_n31; 
@(negedge clk)
!Wreq && !Nreq  &&   Lreq  &&   Lflit_id[2] |->  (nextstate[1]);
endproperty

property property_n32; 
@(negedge clk)
!Ereq && !Nreq  &&   Lreq  &&   Nflit_id[2] |->  (nextstate[1]);
endproperty

property property_n33; 
@(negedge clk)
!Ereq && !Nreq  &&   Lreq  &&   Sflit_id[2] |->  (nextstate[1]);
endproperty

property property_n34; 
@(negedge clk)
!Ereq && !Nreq  &&   Lreq  &&   Wflit_id[2] |->  (nextstate[1]);
endproperty

property property_n35; 
@(negedge clk)
!Ereq && !Nreq  &&   Lreq  &&   Eflit_id[2] |->  (nextstate[1]);
endproperty

property property_n36; 
@(negedge clk)
!Ereq && !Nreq  &&   Lreq  &&   Lflit_id[2] |->  (nextstate[1]);
endproperty

property property_n37; 
@(negedge clk)
 Sflit_id[0] && Sreq  &&   Wreq  &&   !Ereq  &&   Nreq  &&   Lreq  &&   !Nflit_id[1] &&   !Nflit_id[2]  &&   !Sflit_id[1] &&   !Sflit_id[2]  &&   Wflit_id[0]  &&   !Wflit_id[1] &&   !Wflit_id[2]  &&   Eflit_id[0]  &&   !Eflit_id[1] &&   !Eflit_id[2]  &&   Nflit_id[0]  &&   Lflit_id[0]  &&   !Lflit_id[1] &&   !Lflit_id[2]  &&   !rst |->  (!nextstate[1]);
endproperty

property property_n38; 
@(negedge clk)
Sflit_id[0] && Sreq  &&   !Wreq  &&   Nreq  &&   Lreq  &&   !Nflit_id[1] &&   !Nflit_id[2]  &&   !Sflit_id[1] &&   !Sflit_id[2]  &&   Wflit_id[0]  &&   !Wflit_id[1] &&   !Wflit_id[2]  &&   Eflit_id[0]  &&   !Eflit_id[1] &&   !Eflit_id[2]  &&   Nflit_id[0]  &&   Lflit_id[0]  &&   !Lflit_id[1] &&   !Lflit_id[2]  &&   !rst |->  (!nextstate[1]);
endproperty

property property_n39; 
@(negedge clk)
Sflit_id[0] && Sreq  &&   !Nreq  &&   Lreq  &&   !Nflit_id[1] &&   !Nflit_id[2]  &&   !Sflit_id[1] &&   !Sflit_id[2]  &&   Wflit_id[0]  &&   !Wflit_id[1] &&   !Wflit_id[2]  &&   Eflit_id[0]  &&   !Eflit_id[1] &&   !Eflit_id[2]  &&   Nflit_id[0]  &&   Lflit_id[0]  &&   !Lflit_id[1] &&   !Lflit_id[2]  &&   !rst |->  (!nextstate[1]);
endproperty

property property_n40; 
@(negedge clk)
 Sflit_id[0] && !Sreq  &&   !Wreq  &&   Ereq  &&   Nreq  &&   Lreq  &&   !Nflit_id[1] &&   !Nflit_id[2]  &&   !Sflit_id[1] &&   !Sflit_id[2]  &&   Wflit_id[0]  &&   !Wflit_id[1] &&   !Wflit_id[2]  &&   Eflit_id[0]  &&   !Eflit_id[1] &&   !Eflit_id[2]  &&   Nflit_id[0]  &&   Lflit_id[0]  &&   !Lflit_id[1] &&   !Lflit_id[2]  &&   !rst |->  (!nextstate[1]);
endproperty

property property_n41; 
@(negedge clk)
 Sreq && Wreq  &&   !Ereq  &&   Nreq  &&   Lreq  &&   !Nflit_id[1] &&   Nflit_id[2]  &&   !Sflit_id[0]  &&   !Sflit_id[1] &&   Sflit_id[2]  &&   !Wflit_id[0]  &&   !Wflit_id[1] &&   Wflit_id[2]  &&   !Eflit_id[0]  &&   !Eflit_id[1] &&   Eflit_id[2]  &&   !Nflit_id[0]  &&   !Lflit_id[0]  &&   !Lflit_id[1] &&   Lflit_id[2]  &&   !rst |->  (!nextstate[1]);
endproperty

property property_n42; 
@(negedge clk)
Sreq && Wreq  &&   !Ereq  &&   Lreq  &&   !Nflit_id[2]  &&   !Sflit_id[0]  &&   Sflit_id[1] &&   !Sflit_id[2]  &&   !Wflit_id[0]  &&   Wflit_id[1] &&   !Wflit_id[2]  &&   !Eflit_id[0]  &&   Eflit_id[1] &&   !Eflit_id[2]  &&   !Nflit_id[0]  &&   Nflit_id[1] &&   !Lflit_id[0]  &&   Lflit_id[1] &&   !Lflit_id[2]  &&   !rst |->  (!nextstate[1]);
endproperty

property property_n43; 
@(negedge clk)
Sreq && !Wreq  &&   Nreq  &&   Lreq  &&   !Nflit_id[1] &&   Nflit_id[2]  &&   !Sflit_id[0]  &&   !Sflit_id[1] &&   Sflit_id[2]  &&   !Wflit_id[0]  &&   !Wflit_id[1] &&   Wflit_id[2]  &&   !Eflit_id[0]  &&   !Eflit_id[1] &&   Eflit_id[2]  &&   !Nflit_id[0]  &&   !Lflit_id[0]  &&   !Lflit_id[1] &&   Lflit_id[2]  &&   !rst |->  (!nextstate[1]);
endproperty

property property_n44; 
@(negedge clk)
Sreq && Ereq  &&   !Nreq  &&   Lreq  &&   !Nflit_id[1] &&   Nflit_id[2]  &&   !Sflit_id[0]  &&   !Sflit_id[1] &&   Sflit_id[2]  &&   !Wflit_id[0]  &&   !Wflit_id[1] &&   Wflit_id[2]  &&   !Eflit_id[0]  &&   !Eflit_id[1] &&   Eflit_id[2]  &&   !Nflit_id[0]  &&   !Lflit_id[0]  &&   !Lflit_id[1] &&   Lflit_id[2]  &&   !rst |->  (!nextstate[1]);
endproperty

property property_n45; 
@(negedge clk)
!Lreq && !rst |->  (!nextstate[1]);
endproperty

property property_n46; 
@(negedge clk)
rst |-> (!nextstate[1]);
endproperty

property property_n47; 
@(negedge clk)
!Sreq && !Ereq  &&   Nreq  &&   Lflit_id[0]  |->  (nextstate[2]);
endproperty


property property_n48; 
@(negedge clk)
!Wreq && Ereq  &&   Nreq  &&   !Lreq  &&   Nflit_id[2] |->  (nextstate[2]);
endproperty

property property_n49; 
@(negedge clk)
!Wreq && Ereq  &&   Nreq  &&   !Lreq  &&   Sflit_id[2] |->  (nextstate[2]);
endproperty

property property_n50; 
@(negedge clk)
!Wreq && Ereq  &&   Nreq  &&   !Lreq  &&   Wflit_id[2] |->  (nextstate[2]);
endproperty

property property_n51; 
@(negedge clk)
!Wreq && Ereq  &&   Nreq  &&   !Lreq  &&   Eflit_id[2] |->  (nextstate[2]);
endproperty

property property_n52; 
@(negedge clk)
!Wreq && Ereq  &&   Nreq  &&   !Lreq  &&   Lflit_id[2] |->  (nextstate[2]);
endproperty

property property_n53; 
@(negedge clk)
!Ereq && Nreq  &&   !Lreq  &&   Lflit_id[0] |-> (nextstate[2]);
endproperty

property property_n54; 
@(negedge clk)
Sreq && !Wreq  &&   Ereq  &&   Nreq  &&   Lreq  &&   !Nflit_id[2]  &&   !Sflit_id[0]  &&   Sflit_id[1] &&   !Sflit_id[2]  &&   !Wflit_id[0]  &&   Wflit_id[1] &&   !Wflit_id[2]  &&   !Eflit_id[0]  &&   Eflit_id[1] &&   !Eflit_id[2]  &&   !Nflit_id[0]  &&   Nflit_id[1] &&   !Lflit_id[0]  &&   Lflit_id[1] &&   !Lflit_id[2]  &&   !rst |->  (!nextstate[2]);
endproperty

property property_n55; 
@(negedge clk)
!Sreq && Wreq  &&   Ereq  &&   Nreq  &&   Lreq  &&   !Nflit_id[1] &&   Nflit_id[2]  &&   !Sflit_id[0]  &&   !Sflit_id[1] &&   Sflit_id[2]  &&   !Wflit_id[0]  &&   !Wflit_id[1] &&   Wflit_id[2]  &&   !Eflit_id[0]  &&   !Eflit_id[1] &&   Eflit_id[2]  &&   !Nflit_id[0]  &&   !Lflit_id[0]  &&   !Lflit_id[1] &&   Lflit_id[2]  &&   !rst |->  (!nextstate[2]);
endproperty

property property_n56; 
@(negedge clk)
!Sreq && Wreq  &&   Ereq  &&   Nreq  &&   Lreq  &&   !Nflit_id[2]  &&   !Sflit_id[2]  &&   !Wflit_id[2]  &&   !Eflit_id[2]  &&   Lflit_id[1] &&   !Lflit_id[2]  &&   !rst |->  (!nextstate[2]);
endproperty

property property_n57; 
@(negedge clk)
!Sreq && !Wreq  &&   Nreq  &&   Lreq  &&   !Nflit_id[2]  &&   !Sflit_id[0]  &&   Sflit_id[1] &&   !Sflit_id[2]  &&   !Wflit_id[0]  &&   Wflit_id[1] &&   !Wflit_id[2]  &&   !Eflit_id[0]  &&   Eflit_id[1] &&   !Eflit_id[2]  &&   !Nflit_id[0]  &&   Nflit_id[1] &&   !Lflit_id[0]  &&   Lflit_id[1] &&   !Lflit_id[2]  &&   !rst |->  (!nextstate[2]);
endproperty

property property_n58; 
@(negedge clk)
Wreq && !Ereq  &&   Nreq  &&   Lreq  &&   !Nflit_id[1] &&   Nflit_id[2]  &&   !Sflit_id[0]  &&   !Sflit_id[1] &&   Sflit_id[2]  &&   !Wflit_id[0]  &&   !Wflit_id[1] &&   Wflit_id[2]  &&   !Eflit_id[0]  &&   !Eflit_id[1] &&   Eflit_id[2]  &&   !Nflit_id[0]  &&   !Lflit_id[0]  &&   !Lflit_id[1] &&   Lflit_id[2]  &&   !rst |->  (!nextstate[2]);
endproperty

property property_n59; 
@(negedge clk)
!Wreq && Nreq  &&   Lreq  &&   !Sflit_id[0]  &&   !Wflit_id[0]  &&   !Eflit_id[0]  &&   !Nflit_id[0]  &&   !Lflit_id[0]  &&   Lflit_id[2]  &&   !rst |->  (!nextstate[2]);
endproperty

property property_n60; 
@(negedge clk)
!Wreq && Nreq  &&   Lreq  &&   Lflit_id[0]  &&   !rst |->  (!nextstate[2]);
endproperty

property property_n61; 
@(negedge clk)
!Nreq && !rst |->  (!nextstate[2]);
endproperty

property property_n62; 
@(negedge clk)
rst |-> (!nextstate[2]);
endproperty

property property_n63; 
@(negedge clk)
Sflit_id[0] && !Sreq  &&   !Wreq  &&   Ereq  &&   Lreq |->  (nextstate[3]);
endproperty

property property_n64; 
@(negedge clk)
Sflit_id[0] && !Sreq  &&   !Wreq  &&   Nreq  &&   Lreq |->  (nextstate[3]);
endproperty

property property_n65; 
@(negedge clk)
!Sreq && !Wreq  &&   Ereq  &&   Lreq  &&   Wflit_id[0]  |-> (nextstate[3]);
endproperty

property property_n66; 
@(negedge clk)
!Sreq && !Wreq  &&   Ereq  &&   Lreq  &&   Eflit_id[0]  |-> (nextstate[3]);
endproperty

property property_n67; 
@(negedge clk)
!Sreq && !Wreq  &&   Ereq  &&   Lreq  &&   Nflit_id[0] |-> (nextstate[3]);
endproperty

property property_n68; 
@(negedge clk)
!Sreq && !Wreq  &&   Ereq  &&   Lreq  &&   Lflit_id[0] |-> (nextstate[3]);
endproperty

property property_n69; 
@(negedge clk)
!Sreq && !Wreq  &&   Nreq  &&   Lreq  &&   Wflit_id[0] |-> (nextstate[3]);
endproperty

property property_n70; 
@(negedge clk)
!Sreq && !Wreq  &&   Nreq  &&   Lreq  &&   Eflit_id[0] |-> (nextstate[3]);
endproperty


property property_n71; 
@(negedge clk)
!Sreq && !Wreq  &&   Nreq  &&   Lreq  &&   Nflit_id[0] |-> (nextstate[3]);
endproperty
 

property property_n72; 
@(negedge clk)
!Sreq && !Wreq  &&   Nreq  &&   Lreq  &&   Lflit_id[0] |-> (nextstate[3]);
endproperty
 

property property_n73; 
@(negedge clk)
Wreq && !Nreq  &&   Lreq  &&   Nflit_id[2] |->  (nextstate[3]);
endproperty

property property_n74; 
@(negedge clk)
Wreq && !Nreq  &&   Lreq  &&   Sflit_id[2] |->  (nextstate[3]);
endproperty

property property_n75; 
@(negedge clk)
Wreq && !Nreq  &&   Lreq  &&   Wflit_id[2] |->  (nextstate[3]);
endproperty

property property_n76; 
@(negedge clk)
Wreq && !Nreq  &&   Lreq  &&   Eflit_id[2] |->  (nextstate[3]);
endproperty

property property_n77; 
@(negedge clk)
Wreq && !Nreq  &&   Lreq  &&   Lflit_id[2] |->  (nextstate[3]);
endproperty

property property_n78; 
@(negedge clk)
!Wreq && Ereq  &&   !Nreq  &&   Lflit_id[0]  |-> (nextstate[3]);
endproperty


property property_n79; 
@(negedge clk)
!Wreq && Ereq  &&   !Nreq  &&   !Lflit_id[2] |->  (nextstate[3]);
endproperty

property property_n80; 
@(negedge clk)
Ereq && !Nreq  &&   Lreq  &&   Nflit_id[2] |->  (nextstate[3]);
endproperty

property property_n81; 
@(negedge clk)
Ereq && !Nreq  &&   Lreq  &&   Sflit_id[2] |->  (nextstate[3]);
endproperty

property property_n82; 
@(negedge clk)
Ereq && !Nreq  &&   Lreq  &&   Wflit_id[2] |->  (nextstate[3]);
endproperty

property property_n83; 
@(negedge clk)
Ereq && !Nreq  &&   Lreq  &&   Eflit_id[2] |->  (nextstate[3]);
endproperty

property property_n84; 
@(negedge clk)
Ereq && !Nreq  &&   Lreq  &&   Lflit_id[2] |->  (nextstate[3]);
endproperty

property property_n85; 
@(negedge clk)
Sflit_id[0] && Sreq  &&   !Wreq  &&   Ereq  &&   Nreq  &&   Lreq  &&   !Nflit_id[1] &&   !Nflit_id[2]  &&   !Sflit_id[1] &&   !Sflit_id[2]  &&   Wflit_id[0]  &&   !Wflit_id[1] &&   !Wflit_id[2]  &&   Eflit_id[0]  &&   !Eflit_id[1] &&   !Eflit_id[2]  &&   Nflit_id[0]  &&   Lflit_id[0]  &&   !Lflit_id[1] &&   !Lflit_id[2]  &&   !rst |->  (!nextstate[3]);
endproperty

property property_n86; 
@(negedge clk)
 Sflit_id[0] && !Sreq  &&   Wreq  &&   Ereq  &&   Nreq  &&   Lreq  &&   !Nflit_id[1] &&   !Nflit_id[2]  &&   !Sflit_id[1] &&   !Sflit_id[2]  &&   Wflit_id[0]  &&   !Wflit_id[1] &&   !Wflit_id[2]  &&   Eflit_id[0]  &&   !Eflit_id[1] &&   !Eflit_id[2]  &&   Nflit_id[0]  &&   Lflit_id[0]  &&   !Lflit_id[1] &&   !Lflit_id[2]  &&   !rst |->  (!nextstate[3]);
endproperty

property property_n87; 
@(negedge clk)
Sreq && !Wreq  &&   Ereq  &&   Nreq  &&   Lreq  &&   !Nflit_id[1] &&   Nflit_id[2]  &&   !Sflit_id[0]  &&   !Sflit_id[1] &&   Sflit_id[2]  &&   !Wflit_id[0]  &&   !Wflit_id[1] &&   Wflit_id[2]  &&   !Eflit_id[0]  &&   !Eflit_id[1] &&   Eflit_id[2]  &&   !Nflit_id[0]  &&   !Lflit_id[0]  &&   !Lflit_id[1] &&   Lflit_id[2]  &&   !rst |->  (!nextstate[3]);
endproperty

property property_n88; 
@(negedge clk)
Sreq && !Wreq  &&   Ereq  &&   Nreq  &&   Lreq  &&   !Nflit_id[2]  &&   !Sflit_id[0]  &&   Sflit_id[1] &&   !Sflit_id[2]  &&   !Wflit_id[0]  &&   Wflit_id[1] &&   !Wflit_id[2]  &&   !Eflit_id[0]  &&   Eflit_id[1] &&   !Eflit_id[2]  &&   !Nflit_id[0]  &&   Nflit_id[1] &&   !Lflit_id[0]  &&   Lflit_id[1] &&   !Lflit_id[2]  &&   !rst |->  (!nextstate[3]);
endproperty

property property_n89; 
@(negedge clk)
!Sreq && Wreq  &&   Ereq  &&   Nreq  &&   Lreq  &&   !Nflit_id[1] &&   Nflit_id[2]  &&   !Sflit_id[0]  &&   !Sflit_id[1] &&   Sflit_id[2]  &&   !Wflit_id[0]  &&   !Wflit_id[1] &&   Wflit_id[2]  &&   !Eflit_id[0]  &&   !Eflit_id[1] &&   Eflit_id[2]  &&   !Nflit_id[0]  &&   !Lflit_id[0]  &&   !Lflit_id[1] &&   Lflit_id[2]  &&   !rst |->  (!nextstate[3]);
endproperty

property property_n90; 
@(negedge clk)
!Sreq && Wreq  &&   Ereq  &&   Nreq  &&   Lreq  &&   !Nflit_id[2]  &&   !Sflit_id[0]  &&   Sflit_id[1] &&   !Sflit_id[2]  &&   !Wflit_id[0]  &&   Wflit_id[1] &&   !Wflit_id[2]  &&   !Eflit_id[0]  &&   Eflit_id[1] &&   !Eflit_id[2]  &&   !Nflit_id[0]  &&   Nflit_id[1] &&   !Lflit_id[0]  &&   Lflit_id[1] &&   !Lflit_id[2]  &&   !rst |->  (!nextstate[3]);
endproperty

property property_n91; 
@(negedge clk)
!Sreq && Wreq  &&   Ereq  &&   Nreq  &&   !Lreq  &&   !Nflit_id[2]  &&   !Sflit_id[2]  &&   !Wflit_id[2]  &&   !Eflit_id[2]  &&   !Lflit_id[2]  &&   !rst |->  (!nextstate[3]);
endproperty

property property_n92; 
@(negedge clk)
!Sreq && Ereq  &&   Nreq  &&   !Lreq  &&   Lflit_id[2]  &&   !rst |->  (!nextstate[3]);
endproperty

property property_n93; 
@(negedge clk)
!Ereq && !rst |->  (!nextstate[3]);
endproperty

property property_n94; 
@(negedge clk)
 rst |-> (!nextstate[3]);
endproperty

property property_n95; 
@(negedge clk)
Sflit_id[0] && Wreq  &&   !Ereq  &&   !Lreq |->  (nextstate[4]);
endproperty

property property_n96; 
@(negedge clk)
Wreq && !Ereq  &&   Lreq  &&   Nflit_id[2] |->  (nextstate[4]);
endproperty

property property_n97; 
@(negedge clk)
Wreq && !Ereq  &&   Lreq  &&   Sflit_id[2] |->  (nextstate[4]);
endproperty

property property_n98; 
@(negedge clk)
Wreq && !Ereq  &&   Lreq  &&   Wflit_id[2] |->  (nextstate[4]);
endproperty

property property_n99; 
@(negedge clk)
Wreq && !Ereq  &&   Lreq  &&   Eflit_id[2] |->  (nextstate[4]);
endproperty

property property_n100; 
@(negedge clk)
Wreq && !Ereq  &&   Lreq  &&   Lflit_id[2] |->  (nextstate[4]);
endproperty

property property_n101; 
@(negedge clk)
Wreq && !Ereq  &&   !Lreq  &&   Wflit_id[0] |-> (nextstate[4]);
endproperty

property property_n102; 
@(negedge clk)
Wreq && !Ereq  &&   !Lreq  &&   Eflit_id[0]  |-> (nextstate[4]);
endproperty


property property_n103; 
@(negedge clk)
Wreq && !Ereq  &&   !Lreq  &&   Nflit_id[0] |-> (nextstate[4]);
endproperty


property property_n104; 
@(negedge clk)
Wreq && !Ereq  &&   !Lreq  &&   Lflit_id[0]  |-> (nextstate[4]);
endproperty

property property_n105; 
@(negedge clk)
Sflit_id[0] && !Sreq  &&   Wreq  &&   Ereq  &&   Lreq  &&   !Nflit_id[1] &&   !Nflit_id[2]  &&   !Sflit_id[1] &&   !Sflit_id[2]  &&   Wflit_id[0]  &&   !Wflit_id[1] &&   !Wflit_id[2]  &&   Eflit_id[0]  &&   !Eflit_id[1] &&   !Eflit_id[2]  &&   Nflit_id[0]  &&   Lflit_id[0]  &&   !Lflit_id[1] &&   !Lflit_id[2]  &&   !rst |->  (!nextstate[4]);
endproperty

property property_n106; 
@(negedge clk)
 Sreq && Wreq  &&   Ereq  &&   !Nreq  &&   Lreq  &&   !Nflit_id[1] &&   Nflit_id[2]  &&   !Sflit_id[0]  &&   !Sflit_id[1] &&   Sflit_id[2]  &&   !Wflit_id[0]  &&   !Wflit_id[1] &&   Wflit_id[2]  &&   !Eflit_id[0]  &&   !Eflit_id[1] &&   Eflit_id[2]  &&   !Nflit_id[0]  &&   !Lflit_id[0]  &&   !Lflit_id[1] &&   Lflit_id[2]  &&   !rst |->  (!nextstate[4]);
endproperty

property property_n107; 
@(negedge clk)
!Sreq && Wreq  &&   Ereq  &&   Lreq  &&   !Nflit_id[1] &&   Nflit_id[2]  &&   !Sflit_id[0]  &&   !Sflit_id[1] &&   Sflit_id[2]  &&   !Wflit_id[0]  &&   !Wflit_id[1] &&   Wflit_id[2]  &&   !Eflit_id[0]  &&   !Eflit_id[1] &&   Eflit_id[2]  &&   !Nflit_id[0]  &&   !Lflit_id[0]  &&   !Lflit_id[1] &&   Lflit_id[2]  &&   !rst |->  (!nextstate[4]);
endproperty

property property_n108; 
@(negedge clk)
Wreq && Ereq  &&   !Nreq  &&   Lreq  &&   !Nflit_id[2]  &&   !Sflit_id[0]  &&   Sflit_id[1] &&   !Sflit_id[2]  &&   !Wflit_id[0]  &&   Wflit_id[1] &&   !Wflit_id[2]  &&   !Eflit_id[0]  &&   Eflit_id[1] &&   !Eflit_id[2]  &&   !Nflit_id[0]  &&   Nflit_id[1] &&   !Lflit_id[0]  &&   Lflit_id[1] &&   !Lflit_id[2]  &&   !rst |->  (!nextstate[4]);
endproperty

property property_n109; 
@(negedge clk)
!Wreq && !rst |->  (!nextstate[4]);
endproperty

property property_n110; 
@(negedge clk)
rst |-> (!nextstate[4]);
endproperty

property property_n111; 
@(negedge clk)
rst |-> ##1 (nextstate[0]);
endproperty

property property_n112; 
@(negedge clk)
Sreq && Wreq  &&   !Ereq  &&   !Nflit_id[2]  &&   !Sflit_id[2]  &&   !Wflit_id[2]  &&   !Eflit_id[2]  &&   !Lflit_id[2]  &&   !rst |->  ##1 (!nextstate[0]);
endproperty

property property_n113; 
@(negedge clk)
Sreq && !Wreq  &&   !Ereq  &&   Nreq  &&   !Nflit_id[2]  &&   !Sflit_id[2]  &&   !Wflit_id[2]  &&   !Eflit_id[2]  &&   !Lflit_id[2]  &&   !rst |->  ##1 (!nextstate[0]);
endproperty

property property_n114; 
@(negedge clk)
Sreq && !Wreq  &&   !Ereq  &&   !Nreq  &&   Lreq  &&   !Nflit_id[2]  &&   !Sflit_id[2]  &&   !Wflit_id[2]  &&   !Eflit_id[2]  &&   !Lflit_id[2]  &&   !rst |->  ##1 (!nextstate[0]);
endproperty

property property_n115; 
@(negedge clk)
Sreq && !Wreq  &&   !Ereq  &&   !Nreq  &&   !Lreq  &&   !Nflit_id[2]  &&   !Sflit_id[2]  &&   !Wflit_id[2]  &&   !Eflit_id[2]  &&   Lflit_id[1] &&   !Lflit_id[2]  &&   !rst|-> ##1(!nextstate[0]);
endproperty

property property_n116; 
@(negedge clk)
Sreq && Ereq  &&   !Nflit_id[2]  &&   !Sflit_id[2]  &&   !Wflit_id[2]  &&   !Eflit_id[2]  &&   !Lflit_id[2]  &&   !rst |->  ##1 (!nextstate[0]);
endproperty

property property_n117; 
@(negedge clk)
Sreq && Lflit_id[2]  &&   !rst|-> ##1(!nextstate[0]);
endproperty

property property_n118; 
@(negedge clk)
!Sreq && Wreq  &&   Ereq  &&   !Nreq  &&   !Lreq  &&   !Nflit_id[2]  &&   !Sflit_id[0]  &&   Sflit_id[1] &&   !Sflit_id[2]  &&   !Wflit_id[0]  &&   Wflit_id[1] &&   !Wflit_id[2]  &&   !Eflit_id[0]  &&   Eflit_id[1] &&   !Eflit_id[2]  &&   !Nflit_id[0]  &&   Nflit_id[1] &&   !Lflit_id[0]  &&   Lflit_id[1] &&   !Lflit_id[2]  &&   !rst|-> ##1(!nextstate[0]);
endproperty

property property_n119; 
@(negedge clk)
!Sreq && Wreq  &&   !Ereq  &&   !Nreq  &&   !Lreq  &&   Lflit_id[2]  &&   !rst|-> ##1(!nextstate[0]);
endproperty

property property_n120; 
@(negedge clk)
!Sreq && Wreq  &&   Nreq  &&   !rst|-> ##1(!nextstate[0]);
endproperty

property property_n121; 
@(negedge clk)
!Sreq && !Wreq  &&   Ereq  &&   Nreq  &&   Lreq  &&   !Sflit_id[0]  &&   !Wflit_id[0]  &&   !Eflit_id[0]  &&   !Nflit_id[0]  &&   !Lflit_id[0]  &&   !Lflit_id[2]  &&   !rst|-> ##1(!nextstate[0]);
endproperty

property property_n122; 
@(negedge clk)
!Sreq && !Wreq  &&   Ereq  &&   Nreq  &&   !Lreq  &&   !Sflit_id[0]  &&   !Wflit_id[0]  &&   !Eflit_id[0]  &&   !Nflit_id[0]  &&   !Lflit_id[0]  &&   !rst|-> ##1(!nextstate[0]);
endproperty

property property_n123; 
@(negedge clk)
!Sreq && !Wreq  &&   Ereq  &&   Nreq  &&   Lflit_id[0]  &&   !rst|-> ##1(!nextstate[0]);
endproperty

property property_n124; 
@(negedge clk)
!Sreq && !Wreq  &&   !Ereq  &&   !Nreq  &&   Lreq  &&   Lflit_id[0]  &&   !rst|-> ##1(!nextstate[0]);
endproperty

property property_n125; 
@(negedge clk)
!Sreq && Ereq  &&   !Nreq  &&   !Lreq  &&   !Sflit_id[0]  &&   !Wflit_id[0]  &&   !Eflit_id[0]  &&   !Nflit_id[0]  &&   !Lflit_id[0]  &&   Lflit_id[2]  &&   !rst|-> ##1(!nextstate[0]);
endproperty

property property_n126; 
@(negedge clk)
!Sreq && Ereq  &&   !Nreq  &&   !Lreq  &&   Lflit_id[0]  &&   !rst|-> ##1(!nextstate[0]);
endproperty

property property_n127; 
@(negedge clk)
Sflit_id[0] && !Sreq  &&   !Wreq  &&   Lreq|-> ##1(nextstate[1]);
endproperty

property property_n128; 
@(negedge clk)
Sflit_id[0] && !Sreq  &&   !Nreq  &&   Lreq|-> ##1(nextstate[1]);
endproperty

property property_n129; 
@(negedge clk)
Sflit_id[0] && !Wreq  &&   Ereq  &&   Lreq|-> ##1(nextstate[1]);
endproperty

property property_n130; 
@(negedge clk)
 Sreq && !Wreq  &&   Ereq  &&   !Nflit_id[2]  &&   !Lflit_id[1]|-> ##1(nextstate[1]);
endproperty

property property_n131; 
@(negedge clk)
 Sreq && !Wreq  &&   Ereq  &&   !Sflit_id[2]  &&   !Lflit_id[1] |->  ##1(nextstate[1]);
endproperty

property property_n132; 
@(negedge clk)
 Sreq && !Wreq  &&   Ereq  &&   !Wflit_id[2]  &&   !Lflit_id[1] |->  ##1(nextstate[1]);
endproperty

property property_n133; 
@(negedge clk)
 Sreq && !Wreq  &&   Ereq  &&   !Eflit_id[2]  &&   !Lflit_id[1] |->  ##1(nextstate[1]);
endproperty

property property_n134; 
@(negedge clk)
 Sreq && !Wreq  &&   Ereq  &&   !Lflit_id[1] &&   !Lflit_id[2] |->  ##1(nextstate[1]);
endproperty

property property_n135; 
@(negedge clk)
!Sreq && Wreq  &&   Lreq  &&   !Sflit_id[0]  &&   !Lflit_id[2] |->  ##1(nextstate[1]);
endproperty

property property_n136; 
@(negedge clk)
!Sreq && Wreq  &&   Lreq  &&   !Wflit_id[0]  &&   !Lflit_id[2] |->  ##1(nextstate[1]);
endproperty

property property_n137; 
@(negedge clk)
!Sreq && Wreq  &&   Lreq  &&   !Eflit_id[0]  &&   !Lflit_id[2] |->  ##1(nextstate[1]);
endproperty

property property_n138; 
@(negedge clk)
!Sreq && Wreq  &&   Lreq  &&   !Nflit_id[0]  &&   !Lflit_id[2] |->  ##1(nextstate[1]);
endproperty

property property_n139; 
@(negedge clk)
!Sreq && Wreq  &&   Lreq  &&   !Lflit_id[0]  &&   !Lflit_id[2] |->  ##1(nextstate[1]);
endproperty

property property_n140; 
@(negedge clk)
!Sreq && !Wreq  &&   Lreq  &&   Wflit_id[0]  |-> ##1 (nextstate[1]);
endproperty

property property_n141; 
@(negedge clk)
!Sreq && !Wreq  &&   Lreq  &&   Eflit_id[0]  |-> ##1 (nextstate[1]);
endproperty

property property_n142; 
@(negedge clk)
!Sreq && !Wreq  &&   Lreq  &&   Nflit_id[0]  |-> ##1 (nextstate[1]);
endproperty

property property_n143; 
@(negedge clk)
!Sreq && !Wreq  &&   Lreq  &&   Lflit_id[0]  |-> ##1 (nextstate[1]);
endproperty

property property_n144; 
@(negedge clk)
!Sreq && !Nreq  &&   Lreq  &&   Wflit_id[0]  |-> ##1 (nextstate[1]);
endproperty

property property_n145; 
@(negedge clk)
!Sreq && !Nreq  &&   Lreq  &&   Eflit_id[0]  |-> ##1 (nextstate[1]);
endproperty

property property_n146; 
@(negedge clk)
!Sreq && !Nreq  &&   Lreq  &&   Nflit_id[0] |-> ##1 (nextstate[1]);
endproperty

property property_n147; 
@(negedge clk)
!Sreq && !Nreq  &&   Lreq  &&   Lflit_id[0]  |-> ##1 (nextstate[1]);
endproperty



property property_n148; 
@(negedge clk)
!Wreq && Ereq  &&   Lreq  &&   !Nflit_id[2]  &&   !Lflit_id[1] |->  ##1(nextstate[1]);
endproperty

property property_n149; 
@(negedge clk)
!Wreq && Ereq  &&   Lreq  &&   !Sflit_id[2]  &&   !Lflit_id[1] |->  ##1(nextstate[1]);
endproperty

property property_n150; 
@(negedge clk)
!Wreq && Ereq  &&   Lreq  &&   Wflit_id[0] |-> ##1 (nextstate[1]);
endproperty

property property_n151; 
@(negedge clk)
!Wreq && Ereq  &&   Lreq  &&   !Wflit_id[2]  &&   !Lflit_id[1] |->  ##1(nextstate[1]);
endproperty

property property_n152; 
@(negedge clk)
!Wreq && Ereq  &&   Lreq  &&   Eflit_id[0]  |-> ##1 (nextstate[1]);
endproperty

property property_n153; 
@(negedge clk)
!Wreq && Ereq  &&   Lreq  &&   !Eflit_id[2]  &&   !Lflit_id[1]|-> ##1(nextstate[1]);
endproperty

property property_n154; 
@(negedge clk)
!Wreq && Ereq  &&   Lreq  &&   Nflit_id[0]  |-> ##1 (nextstate[1]);
endproperty

property property_n155; 
@(negedge clk)
!Wreq && Ereq  &&   Lreq  &&   Lflit_id[0]  |-> ##1 (nextstate[1]);
endproperty

property property_n156; 
@(negedge clk)
!Wreq && Ereq  &&   Lreq  &&   !Lflit_id[1] &&   !Lflit_id[2] |->  ##1(nextstate[1]);
endproperty

property property_n157; 
@(negedge clk)
Sreq && Wreq  &&   !Ereq  &&   Lreq  &&   !Nflit_id[2]  &&   !Sflit_id[0]  &&   Sflit_id[1] &&   !Sflit_id[2]  &&   !Wflit_id[0]  &&   Wflit_id[1] &&   !Wflit_id[2]  &&   !Eflit_id[0]  &&   Eflit_id[1] &&   !Eflit_id[2]  &&   !Nflit_id[0]  &&   Nflit_id[1] &&   !Lflit_id[0]  &&   Lflit_id[1] &&   !Lflit_id[2]  &&   !rst|-> ##1(!nextstate[1]);
endproperty

property property_n158; 
@(negedge clk)
Sreq && !Wreq  &&   Ereq  &&   Nreq  &&   Lreq  &&   !Nflit_id[1] &&   Nflit_id[2]  &&   !Sflit_id[0]  &&   !Sflit_id[1] &&   Sflit_id[2]  &&   !Wflit_id[0]  &&   !Wflit_id[1] &&   Wflit_id[2]  &&   !Eflit_id[0]  &&   !Eflit_id[1] &&   Eflit_id[2]  &&   !Nflit_id[0]  &&   !Lflit_id[0]  &&   !Lflit_id[1] &&   Lflit_id[2]  &&   !rst|-> ##1(!nextstate[1]);
endproperty

property property_n159; 
@(negedge clk)
Sreq && Ereq  &&   !Nreq  &&   Lreq  &&   !Nflit_id[2]  &&   !Sflit_id[2]  &&   !Wflit_id[2]  &&   !Eflit_id[2]  &&   !Lflit_id[2]  &&   !rst|-> ##1(!nextstate[1]);
endproperty

property property_n160; 
@(negedge clk)
Sreq && !Ereq  &&   Nreq  &&   Lreq  &&   !Nflit_id[1] &&   Nflit_id[2]  &&   !Sflit_id[0]  &&   !Sflit_id[1] &&   Sflit_id[2]  &&   !Wflit_id[0]  &&   !Wflit_id[1] &&   Wflit_id[2]  &&   !Eflit_id[0]  &&   !Eflit_id[1] &&   Eflit_id[2]  &&   !Nflit_id[0]  &&   !Lflit_id[0]  &&   !Lflit_id[1] &&   Lflit_id[2]  &&   !rst|-> ##1(!nextstate[1]);
endproperty

property property_n161; 
@(negedge clk)
Sreq && !Ereq  &&   Lreq  &&   !Nflit_id[2]  &&   !Sflit_id[2]  &&   !Wflit_id[2]  &&   !Eflit_id[2]  &&   !Lflit_id[1] &&   !Lflit_id[2]  &&   !rst|-> ##1(!nextstate[1]);
endproperty

property property_n162; 
@(negedge clk)
Sreq && !Nreq  &&   Lreq  &&   !Nflit_id[1] &&   Nflit_id[2]  &&   !Sflit_id[0]  &&   !Sflit_id[1] &&   Sflit_id[2]  &&   !Wflit_id[0]  &&   !Wflit_id[1] &&   Wflit_id[2]  &&   !Eflit_id[0]  &&   !Eflit_id[1] &&   Eflit_id[2]  &&   !Nflit_id[0]  &&   !Lflit_id[0]  &&   !Lflit_id[1] &&   Lflit_id[2]  &&   !rst|-> ##1(!nextstate[1]);
endproperty

property property_n163; 
@(negedge clk)
Sreq && !Lreq  &&   !rst|-> ##1(!nextstate[1]);
endproperty

property property_n164; 
@(negedge clk)
!Sreq && Wreq  &&   !Lreq  &&   !Sflit_id[0]  &&   !Wflit_id[0]  &&   !Eflit_id[0]  &&   !Nflit_id[0]  &&   !Lflit_id[0]  &&   !rst|-> ##1(!nextstate[1]);
endproperty

property property_n165; 
@(negedge clk)
!Sreq && !Wreq  &&   Ereq  &&   !Nreq  &&   !Lreq  &&   !Sflit_id[0]  &&   !Wflit_id[0]  &&   !Eflit_id[0]  &&   !Nflit_id[0]  &&   !Lflit_id[0]  &&   !rst|-> ##1(!nextstate[1]);
endproperty

property property_n166; 
@(negedge clk)
!Sreq && !Wreq  &&   !Ereq  &&   Nreq  &&   !Lreq  &&   !Nflit_id[2]  &&   !Sflit_id[0]  &&   Sflit_id[1] &&   !Sflit_id[2]  &&   !Wflit_id[0]  &&   Wflit_id[1] &&   !Wflit_id[2]  &&   !Eflit_id[0]  &&   Eflit_id[1] &&   !Eflit_id[2]  &&   !Nflit_id[0]  &&   Nflit_id[1] &&   !Lflit_id[0]  &&   Lflit_id[1] &&   !Lflit_id[2]  &&   !rst|-> ##1(!nextstate[1]);
endproperty

property property_n167; 
@(negedge clk)
!Sreq && !Wreq  &&   Nreq  &&   Lreq  &&   !Sflit_id[0]  &&   !Wflit_id[0]  &&   !Eflit_id[0]  &&   !Nflit_id[0]  &&   !Lflit_id[0]  &&   Lflit_id[2]  &&   !rst|-> ##1(!nextstate[1]);
endproperty

property property_n168; 
@(negedge clk)
!Sreq && !Wreq  &&   Nreq  &&   !Lreq  &&   !Sflit_id[0]  &&   !Wflit_id[0]  &&   !Eflit_id[0]  &&   !Nflit_id[0]  &&   !Lflit_id[0]  &&   Lflit_id[2]  &&   !rst|-> ##1(!nextstate[1]);
endproperty

property property_n169; 
@(negedge clk)
!Sreq && !Lreq  &&   Lflit_id[0]  &&   !rst|-> ##1(!nextstate[1]);
endproperty

property property_n170; 
@(negedge clk)
 rst |-> ##1 (!nextstate[1]);
endproperty

property property_n171; 
@(negedge clk)
Sflit_id[0] && Wreq  &&   Nreq  &&   !Lreq|-> ##1(nextstate[2]);
endproperty

property property_n172; 
@(negedge clk)
Sflit_id[0] && Ereq  &&   Nreq  &&   !Lreq|-> ##1(nextstate[2]);
endproperty

property property_n173; 
@(negedge clk)
Wreq && Nreq  &&   !Lreq  &&   Wflit_id[0]|->  ##1 (nextstate[2]);
endproperty

property property_n174; 
@(negedge clk)
Wreq && Nreq  &&   !Lreq  &&   Eflit_id[0]  |-> ##1 (nextstate[2]);
endproperty

property property_n175; 
@(negedge clk)
Wreq && Nreq  &&   !Lreq  &&   Nflit_id[0]  |-> ##1 (nextstate[2]);
endproperty

property property_n176; 
@(negedge clk)
Wreq && Nreq  &&   !Lreq  &&   Lflit_id[0]  |-> ##1 (nextstate[2]);
endproperty

property property_n177; 
@(negedge clk)
!Wreq && Ereq  &&   Nreq  &&   !Lreq  &&   !Nflit_id[1] |-> ##1(nextstate[2]);
endproperty

property property_n178; 
@(negedge clk)
!Wreq && Ereq  &&   Nreq  &&   !Lreq  &&   Nflit_id[2] |-> ##1(nextstate[2]);
endproperty

property property_n179; 
@(negedge clk)
!Wreq && Ereq  &&   Nreq  &&   !Lreq  &&   !Sflit_id[1] |-> ##1(nextstate[2]);
endproperty

property property_n180; 
@(negedge clk)
!Wreq && Ereq  &&   Nreq  &&   !Lreq  &&   Sflit_id[2] |-> ##1(nextstate[2]);
endproperty

property property_n181; 
@(negedge clk)
!Wreq && Ereq  &&   Nreq  &&   !Lreq  &&   !Wflit_id[1] |->  ##1(nextstate[2]);
endproperty

property property_n182; 
@(negedge clk)
!Wreq && Ereq  &&   Nreq  &&   !Lreq  &&   Wflit_id[2] |->  ##1(nextstate[2]);
endproperty

property property_n183; 
@(negedge clk)
!Wreq && Ereq  &&   Nreq  &&   !Lreq  &&   !Eflit_id[1] |->  ##1(nextstate[2]);
endproperty

property property_n184; 
@(negedge clk)
!Wreq && Ereq  &&   Nreq  &&   !Lreq  &&   Eflit_id[2] |->  ##1(nextstate[2]);
endproperty

property property_n185; 
@(negedge clk)
!Wreq && Ereq  &&   Nreq  &&   !Lreq  &&   !Lflit_id[1] |->  ##1(nextstate[2]);
endproperty

property property_n186; 
@(negedge clk)
!Wreq && Ereq  &&   Nreq  &&   !Lreq  &&   Lflit_id[2] |->  ##1(nextstate[2]);
endproperty

property property_n187; 
@(negedge clk)
Ereq && Nreq  &&   !Lreq  &&   Wflit_id[0]|->  ##1 (nextstate[2]);
endproperty

property property_n188; 
@(negedge clk)
Ereq && Nreq  &&   !Lreq  &&   Eflit_id[0]|->  ##1 (nextstate[2]);
endproperty

property property_n189; 
@(negedge clk)
Ereq && Nreq  &&   !Lreq  &&   Nflit_id[0]|->  ##1 (nextstate[2]);
endproperty

property property_n190; 
@(negedge clk)
Ereq && Nreq  &&   !Lreq  &&   Lflit_id[0]|->  ##1 (nextstate[2]);
endproperty

property property_n191; 
@(negedge clk)
 Sreq && Wreq  &&   !Ereq  &&   Nreq  &&   Lreq  &&   !Nflit_id[1] &&   Nflit_id[2]  &&   !Sflit_id[0]  &&   !Sflit_id[1] &&   Sflit_id[2]  &&   !Wflit_id[0]  &&   !Wflit_id[1] &&   Wflit_id[2]  &&   !Eflit_id[0]  &&   !Eflit_id[1] &&   Eflit_id[2]  &&   !Nflit_id[0]  &&   !Lflit_id[0]  &&   !Lflit_id[1] &&   Lflit_id[2]  &&   !rst|-> ##1(!nextstate[2]);
endproperty

property property_n192; 
@(negedge clk)
 Sreq && !Wreq  &&   !Ereq  &&   Nreq  &&   Lreq  &&   !Nflit_id[2]  &&   !Sflit_id[0]  &&   Sflit_id[1] &&   !Sflit_id[2]  &&   !Wflit_id[0]  &&   Wflit_id[1] &&   !Wflit_id[2]  &&   !Eflit_id[0]  &&   Eflit_id[1] &&   !Eflit_id[2]  &&   !Nflit_id[0]  &&   Nflit_id[1] &&   !Lflit_id[0]  &&   Lflit_id[1] &&   !Lflit_id[2]  &&   !rst|-> ##1(!nextstate[2]);
endproperty

property property_n193; 
@(negedge clk)
Sreq && !Nreq  &&   !Nflit_id[2]  &&   !Sflit_id[2]  &&   !Wflit_id[2]  &&   !Eflit_id[2]  &&   !Lflit_id[2]  &&   !rst|-> ##1(!nextstate[2]);
endproperty

property property_n194; 
@(negedge clk)
!Sreq && Wreq  &&   Ereq  &&   Nreq  &&   Lreq  &&   !Sflit_id[0]  &&   !Wflit_id[0]  &&   !Eflit_id[0]  &&   !Nflit_id[0]  &&   !Lflit_id[0]  &&   !Lflit_id[2]  &&   !rst|-> ##1(!nextstate[2]);
endproperty

property property_n195; 
@(negedge clk)
!Sreq && Wreq  &&   Ereq  &&   Nreq  &&   Lreq  &&   Lflit_id[0]  &&   !rst|-> ##1(!nextstate[2]);
endproperty

property property_n196; 
@(negedge clk)
!Sreq && Wreq  &&   !Ereq  &&   !Nreq  &&   !Lreq  &&   !Nflit_id[2]  &&   !Sflit_id[0]  &&   Sflit_id[1] &&   !Sflit_id[2]  &&   !Wflit_id[0]  &&   Wflit_id[1] &&   !Wflit_id[2]  &&   !Eflit_id[0]  &&   Eflit_id[1] &&   !Eflit_id[2]  &&   !Nflit_id[0]  &&   Nflit_id[1] &&   !Lflit_id[0]  &&   Lflit_id[1] &&   !Lflit_id[2]  &&   !rst|-> ##1(!nextstate[2]);
endproperty

property property_n197; 
@(negedge clk)
!Sreq && !Wreq  &&   Nreq  &&   Lreq  &&   !Nflit_id[2]  &&   !Sflit_id[0]  &&   Sflit_id[1] &&   !Sflit_id[2]  &&   !Wflit_id[0]  &&   Wflit_id[1] &&   !Wflit_id[2]  &&   !Eflit_id[0]  &&   Eflit_id[1] &&   !Eflit_id[2]  &&   !Nflit_id[0]  &&   Nflit_id[1] &&   !Lflit_id[0]  &&   Lflit_id[1] &&   !Lflit_id[2]  &&   !rst|-> ##1(!nextstate[2]);
endproperty

property property_n198; 
@(negedge clk)
!Sreq && Ereq  &&   !Nreq  &&   !Nflit_id[2]  &&   !Sflit_id[2]  &&   !Wflit_id[2]  &&   !Eflit_id[2]  &&   !Lflit_id[2]  &&   !rst|-> ##1(!nextstate[2]);
endproperty

property property_n199; 
@(negedge clk)
!Sreq && !Ereq  &&   !Nreq  &&   Lreq  &&   !Nflit_id[2]  &&   !Sflit_id[0]  &&   Sflit_id[1] &&   !Sflit_id[2]  &&   !Wflit_id[0]  &&   Wflit_id[1] &&   !Wflit_id[2]  &&   !Eflit_id[0]  &&   Eflit_id[1] &&   !Eflit_id[2]  &&   !Nflit_id[0]  &&   Nflit_id[1] &&   !Lflit_id[0]  &&   Lflit_id[1] &&   !Lflit_id[2]  &&   !rst|-> ##1(!nextstate[2]);
endproperty

property property_n200; 
@(negedge clk)
!Sreq && !Ereq  &&   !Nreq  &&   !Nflit_id[2]  &&   !Sflit_id[2]  &&   !Wflit_id[2]  &&   !Eflit_id[2]  &&   !Lflit_id[1] &&   !Lflit_id[2]  &&   !rst|-> ##1(!nextstate[2]);
endproperty

property property_n201; 
@(negedge clk)
!Wreq && Nreq  &&   Lreq  &&   !Sflit_id[0]  &&   !Wflit_id[0]  &&   !Eflit_id[0]  &&   !Nflit_id[0]  &&   !Lflit_id[0]  &&   Lflit_id[2]  &&   !rst|-> ##1(!nextstate[2]);
endproperty

property property_n202; 
@(negedge clk)
!Wreq && Nreq  &&   Lreq  &&   Lflit_id[0]  &&   !rst|-> ##1(!nextstate[2]);
endproperty

property property_n203; 
@(negedge clk)
!Nreq && Lflit_id[2]  &&   !rst|-> ##1(!nextstate[2]);
endproperty

property property_n204; 
@(negedge clk)
 rst |-> ##1 (!nextstate[2]);
endproperty

property property_n205; 
@(negedge clk)
Wreq && !Nreq  &&   Lreq  &&   Sflit_id[1] |->  ##1(nextstate[3]);
endproperty

property property_n206; 
@(negedge clk)
Wreq && !Nreq  &&   Lreq  &&   Wflit_id[1] |->  ##1(nextstate[3]);
endproperty

property property_n207; 
@(negedge clk)
Wreq && !Nreq  &&   Lreq  &&   Eflit_id[1] |->  ##1(nextstate[3]);
endproperty

property property_n208; 
@(negedge clk)
Wreq && !Nreq  &&   Lreq  &&   Nflit_id[1] |->  ##1(nextstate[3]);
endproperty

property property_n209; 
@(negedge clk)
Wreq && !Nreq  &&   Lreq  &&   Lflit_id[1] |->  ##1(nextstate[3]);
endproperty

property property_n210; 
@(negedge clk)
!Wreq && Ereq  &&   !Nreq  &&   Lflit_id[0]  |-> ##1 (nextstate[3]) ;
endproperty
 

property property_n211; 
@(negedge clk)
!Wreq && Ereq  &&   !Nreq  &&   Lflit_id[2] |->  ##1(nextstate[3]);
endproperty

property property_n212; 
@(negedge clk)
Ereq && !Nreq  &&   Lreq  &&   Sflit_id[1] |->  ##1(nextstate[3]);
endproperty

property property_n213; 
@(negedge clk)
Ereq && !Nreq  &&   Lreq  &&   Wflit_id[1] |->  ##1(nextstate[3]);
endproperty

property property_n214; 
@(negedge clk)
Ereq && !Nreq  &&   Lreq  &&   Eflit_id[1] |->  ##1(nextstate[3]);
endproperty

property property_n215; 
@(negedge clk)
Ereq && !Nreq  &&   Lreq  &&   Nflit_id[1] |->  ##1(nextstate[3]);
endproperty

property property_n216; 
@(negedge clk)
Ereq && !Nreq  &&   Lreq  &&   Lflit_id[1] |->  ##1(nextstate[3]);
endproperty

property property_n217; 
@(negedge clk)
Sreq && !Wreq  &&   Ereq  &&   Nreq  &&   Lreq  &&   !Nflit_id[1] &&   !Sflit_id[1] &&   !Wflit_id[1] &&   !Eflit_id[1] &&   !Lflit_id[1] &&   !rst|-> ##1(!nextstate[3]);
endproperty

property property_n218; 
@(negedge clk)
 Sreq && !Wreq  &&   Ereq  &&   Nreq  &&   Lreq  &&   !Nflit_id[2]  &&   !Sflit_id[0]  &&   Sflit_id[1] &&   !Sflit_id[2]  &&   !Wflit_id[0]  &&   Wflit_id[1] &&   !Wflit_id[2]  &&   !Eflit_id[0]  &&   Eflit_id[1] &&   !Eflit_id[2]  &&   !Nflit_id[0]  &&   Nflit_id[1] &&   !Lflit_id[0]  &&   Lflit_id[1] &&   !Lflit_id[2]  &&   !rst|-> ##1(!nextstate[3]);
endproperty

property property_n219; 
@(negedge clk)
 Sreq && !Wreq  &&   !Ereq  &&   !Nreq  &&   Lreq  &&   !Nflit_id[2]  &&   !Sflit_id[0]  &&   Sflit_id[1] &&   !Sflit_id[2]  &&   !Wflit_id[0]  &&   Wflit_id[1] &&   !Wflit_id[2]  &&   !Eflit_id[0]  &&   Eflit_id[1] &&   !Eflit_id[2]  &&   !Nflit_id[0]  &&   Nflit_id[1] &&   !Lflit_id[0]  &&   Lflit_id[1] &&   !Lflit_id[2]  &&   !rst|-> ##1(!nextstate[3]);
endproperty

property property_n220; 
@(negedge clk)
Sreq && !Wreq  &&   !Ereq  &&   !Lreq  &&   !Nflit_id[2]  &&   !Sflit_id[2]  &&   !Wflit_id[2]  &&   !Eflit_id[2]  &&   !Lflit_id[2]  &&   !rst|-> ##1(!nextstate[3]);
endproperty

property property_n221; 
@(negedge clk)
!Sreq && Wreq  &&   Ereq  &&   Nreq  &&   Lreq  &&   !Nflit_id[1] &&   Nflit_id[2]  &&   !Sflit_id[0]  &&   !Sflit_id[1] &&   Sflit_id[2]  &&   !Wflit_id[0]  &&   !Wflit_id[1] &&   Wflit_id[2]  &&   !Eflit_id[0]  &&   !Eflit_id[1] &&   Eflit_id[2]  &&   !Nflit_id[0]  &&   !Lflit_id[0]  &&   !Lflit_id[1] &&   Lflit_id[2]  &&   !rst|-> ##1(!nextstate[3]);
endproperty

property property_n222; 
@(negedge clk)
!Sreq && Wreq  &&   Ereq  &&   Nreq  &&   Lreq  &&   !Nflit_id[2]  &&   !Sflit_id[0]  &&   Sflit_id[1] &&   !Sflit_id[2]  &&   !Wflit_id[0]  &&   Wflit_id[1] &&   !Wflit_id[2]  &&   !Eflit_id[0]  &&   Eflit_id[1] &&   !Eflit_id[2]  &&   !Nflit_id[0]  &&   Nflit_id[1] &&   !Lflit_id[0]  &&   Lflit_id[1] &&   !Lflit_id[2]  &&   !rst|-> ##1(!nextstate[3]);
endproperty

property property_n223; 
@(negedge clk)
!Sreq && Wreq  &&   Ereq  &&   Nreq  &&   !Lreq  &&   !Nflit_id[2]  &&   !Sflit_id[0]  &&   Sflit_id[1] &&   !Sflit_id[2]  &&   !Wflit_id[0]  &&   Wflit_id[1] &&   !Wflit_id[2]  &&   !Eflit_id[0]  &&   Eflit_id[1] &&   !Eflit_id[2]  &&   !Nflit_id[0]  &&   Nflit_id[1] &&   !Lflit_id[0]  &&   Lflit_id[1] &&   !Lflit_id[2]  &&   !rst|-> ##1(!nextstate[3]);
endproperty

property property_n224; 
@(negedge clk)
!Sreq && !Wreq  &&   !Ereq  &&   Nreq  &&   !Lreq  &&   !Nflit_id[2]  &&   !Sflit_id[2]  &&   !Wflit_id[2]  &&   !Eflit_id[2]  &&   !Lflit_id[2]  &&   !rst|-> ##1(!nextstate[3]);
endproperty

property property_n225; 
@(negedge clk)
!Sreq && !Wreq  &&   !Ereq  &&   !Nreq  &&   !Lreq  &&   !Nflit_id[2]  &&   !Sflit_id[2]  &&   !Wflit_id[2]  &&   !Eflit_id[2]  &&   Lflit_id[1] &&   !Lflit_id[2]  &&   !rst|-> ##1(!nextstate[3]);
endproperty

property property_n226; 
@(negedge clk)
!Sreq && !Wreq  &&   !Ereq  &&   Lreq  &&   !Nflit_id[2]  &&   !Sflit_id[0]  &&   Sflit_id[1] &&   !Sflit_id[2]  &&   !Wflit_id[0]  &&   Wflit_id[1] &&   !Wflit_id[2]  &&   !Eflit_id[0]  &&   Eflit_id[1] &&   !Eflit_id[2]  &&   !Nflit_id[0]  &&   Nflit_id[1] &&   !Lflit_id[0]  &&   Lflit_id[1] &&   !Lflit_id[2]  &&   !rst|-> ##1(!nextstate[3]);
endproperty

property property_n227; 
@(negedge clk)
!Sreq && Ereq  &&   Nreq  &&   Lreq  &&   !Nflit_id[1] &&   !Sflit_id[1] &&   !Wflit_id[1] &&   !Eflit_id[1] &&   !Lflit_id[1] &&   !Lflit_id[2]  &&   !rst|-> ##1(!nextstate[3]);
endproperty

property property_n228; 
@(negedge clk)
!Sreq && Ereq  &&   Nreq  &&   !Lreq  &&   !Nflit_id[2]  &&   !Sflit_id[2]  &&   !Wflit_id[2]  &&   !Eflit_id[2]  &&   !Lflit_id[1] &&   !Lflit_id[2]  &&   !rst|-> ##1(!nextstate[3]);
endproperty

property property_n229; 
@(negedge clk)
!Sreq && Ereq  &&   Nreq  &&   !Lreq  &&   Lflit_id[2]  &&   !rst|-> ##1(!nextstate[3]);
endproperty

property property_n230; 
@(negedge clk)
Wreq && !Ereq  &&   !Nflit_id[2]  &&   !Sflit_id[2]  &&   !Wflit_id[2]  &&   !Eflit_id[2]  &&   !Lflit_id[2]  &&   !rst|-> ##1(!nextstate[3]);
endproperty

property property_n231; 
@(negedge clk)
!Wreq && !Ereq  &&   Lreq  &&   !Nflit_id[2]  &&   !Sflit_id[2]  &&   !Wflit_id[2]  &&   !Eflit_id[2]  &&   !Lflit_id[1] &&   !Lflit_id[2]  &&   !rst|-> ##1(!nextstate[3]);
endproperty

property property_n232; 
@(negedge clk)
!Ereq && Lflit_id[2]  &&   !rst|-> ##1(!nextstate[3]);
endproperty

property property_n233; 
@(negedge clk)
 rst |-> ##1 (!nextstate[3]);
endproperty

property property_n234; 
@(negedge clk)
Wreq && !Ereq  &&   Lflit_id[2] |->  ##1(nextstate[4]);
endproperty

property property_n235; 
@(negedge clk)
 Sflit_id[0] && Sreq  &&   Wreq  &&   Ereq  &&   !Nreq  &&   Lreq  &&   !Nflit_id[1] &&   !Nflit_id[2]  &&   !Sflit_id[1] &&   !Sflit_id[2]  &&   Wflit_id[0]  &&   !Wflit_id[1] &&   !Wflit_id[2]  &&   Eflit_id[0]  &&   !Eflit_id[1] &&   !Eflit_id[2]  &&   Nflit_id[0]  &&   Lflit_id[0]  &&   !Lflit_id[1] &&   !Lflit_id[2]  &&   !rst|-> ##1(!nextstate[4]);
endproperty

property property_n236; 
@(negedge clk)
 Sflit_id[0] && !Sreq  &&   Wreq  &&   Ereq  &&   Nreq  &&   !Lreq  &&   !Nflit_id[1] &&   !Nflit_id[2]  &&   !Sflit_id[1] &&   !Sflit_id[2]  &&   Wflit_id[0]  &&   !Wflit_id[1] &&   !Wflit_id[2]  &&   Eflit_id[0]  &&   !Eflit_id[1] &&   !Eflit_id[2]  &&   Nflit_id[0]  &&   Lflit_id[0]  &&   !Lflit_id[1] &&   !Lflit_id[2]  &&   !rst|-> ##1(!nextstate[4]);
endproperty

property property_n237; 
@(negedge clk)
Sreq && Wreq  &&   Ereq  &&   !Nreq  &&   Lreq  &&   !Sflit_id[0]  &&   !Wflit_id[0]  &&   !Eflit_id[0]  &&   !Nflit_id[0]  &&   !Lflit_id[0]  &&   !Lflit_id[2]  &&   !rst|-> ##1(!nextstate[4]);
endproperty

property property_n238; 
@(negedge clk)
!Sreq && Wreq  &&   Ereq  &&   Lreq  &&   !Sflit_id[0]  &&   !Wflit_id[0]  &&   !Eflit_id[0]  &&   !Nflit_id[0]  &&   !Lflit_id[0]  &&   !rst|-> ##1(!nextstate[4]);
endproperty

property property_n239; 
@(negedge clk)
!Wreq && Ereq  &&   !Nflit_id[2]  &&   !Sflit_id[0]  &&   Sflit_id[1] &&   !Sflit_id[2]  &&   !Wflit_id[0]  &&   Wflit_id[1] &&   !Wflit_id[2]  &&   !Eflit_id[0]  &&   Eflit_id[1] &&   !Eflit_id[2]  &&   !Nflit_id[0]  &&   Nflit_id[1] &&   !Lflit_id[0]  &&   Lflit_id[1] &&   !Lflit_id[2]  &&   !rst|-> ##1(!nextstate[4]);
endproperty

property property_n240; 
@(negedge clk)
!Wreq && !Ereq  &&   Nreq  &&   !Nflit_id[2]  &&   !Sflit_id[0]  &&   Sflit_id[1] &&   !Sflit_id[2]  &&   !Wflit_id[0]  &&   Wflit_id[1] &&   !Wflit_id[2]  &&   !Eflit_id[0]  &&   Eflit_id[1] &&   !Eflit_id[2]  &&   !Nflit_id[0]  &&   Nflit_id[1] &&   !Lflit_id[0]  &&   Lflit_id[1] &&   !Lflit_id[2]  &&   !rst|-> ##1(!nextstate[4]);
endproperty

property property_n241; 
@(negedge clk)
!Wreq && !Ereq  &&   !Nreq  &&   Lreq  &&   !Nflit_id[2]  &&   !Sflit_id[0]  &&   Sflit_id[1] &&   !Sflit_id[2]  &&   !Wflit_id[0]  &&   Wflit_id[1] &&   !Wflit_id[2]  &&   !Eflit_id[0]  &&   Eflit_id[1] &&   !Eflit_id[2]  &&   !Nflit_id[0]  &&   Nflit_id[1] &&   !Lflit_id[0]  &&   Lflit_id[1] &&   !Lflit_id[2]  &&   !rst|-> ##1(!nextstate[4]);
endproperty

property property_n242; 
@(negedge clk)
!Wreq && !Nflit_id[2]  &&   !Sflit_id[2]  &&   !Wflit_id[2]  &&   !Eflit_id[2]  &&   !Lflit_id[1] &&   !Lflit_id[2]  &&   !rst |-> ##1(!nextstate[4]);
endproperty

property property_n243; 
@(negedge clk)
!Wreq && Lflit_id[2]  &&   !rst|-> ##1(!nextstate[4]);
endproperty

property property_n244; 
@(negedge clk)
 rst |-> ##1 (!nextstate[4]);
endproperty


property property_n248; 
@(negedge clk)
!Lflit_id[2] && !Lflit_id[1] &&   !Nflit_id[2]  &&   !Eflit_id[2]  &&   !Wflit_id[2]  &&   !Sflit_id[2]  &&   !Lreq  &&   !Nreq  &&   !Sreq  &&   !rst  &&   Ereq   ##1 !Lflit_id[0] && !Nflit_id[0]  &&   !Eflit_id[0]  &&   !Wflit_id[0]  &&   !Sflit_id[0]  &&   !Lreq  &&   !Nreq  &&   !Sreq  &&   !rst  &&   Ereq |-> ##1(!nextstate[0]);
endproperty

property property_n249; 
@(negedge clk)
!Lflit_id[2] && !Nflit_id[2]  &&   !Eflit_id[2]  &&   !Wflit_id[2]  &&   !Sflit_id[2]  &&   !Lreq  &&   !Wreq  &&   !Sreq  &&   !rst  &&   Nreq  &&   Ereq   ##1 !Lflit_id[0] && !Nflit_id[0]  &&   !Eflit_id[0]  &&   !Wflit_id[0]  &&   !Sflit_id[0]  &&   !Lreq  &&   !Wreq  &&   !Sreq  &&   !rst  &&   Nreq|-> ##1(!nextstate[0]);
endproperty

property property_n251; 
@(negedge clk)
!Lflit_id[2] && !Nflit_id[2]  &&   !Eflit_id[2]  &&   !Wflit_id[2]  &&   !Sflit_id[2]  &&   !Sreq  &&   !rst  &&   Nreq  &&   Wreq   ##1 !Lflit_id[0] && !Nflit_id[0]  &&   !Eflit_id[0]  &&   !Wflit_id[0]  &&   !Sflit_id[0]  &&   !Sreq  &&   !rst  &&   Nreq |-> ##1(!nextstate[0]);
endproperty

property property_n252; 
@(negedge clk)
!Lflit_id[2] && !Nflit_id[2]  &&   !Eflit_id[2]  &&   !Wflit_id[2]  &&   !Sflit_id[2]  &&   !rst  &&   Sreq   ##1 !Lflit_id[0] && !Nflit_id[0]  &&   !Eflit_id[0]  &&   !Wflit_id[0]  &&   !Sflit_id[0]  &&   !rst  &&   Lflit_id[2]  &&   Sreq |-> ##1(!nextstate[0]);
endproperty

property property_n256; 
@(negedge clk)
!Lreq && !Nreq  &&   !Ereq  &&   !rst  &&   Sreq   ##1 !Lreq && !Nreq  &&   !Ereq  &&   !Sreq  &&   !rst  &&   Wreq|-> ##1(!nextstate[0]);
endproperty


property property_n258; 
@(negedge clk)
!Lreq && !Nreq  &&   !Sreq  &&   !rst  &&   Lflit_id[2]  &&   Ereq   ##1 !Lreq && !Nreq  &&   !Sreq  &&   !rst  &&   Ereq|-> ##1 (!nextstate[0]);
endproperty

property property_n260; 
@(negedge clk)
!rst && Lreq   ##1 !Lreq && !Nreq  &&   !Ereq  &&   !Sreq  &&   !rst  &&   Wreq|-> ##1(!nextstate[0]);
endproperty

property property_n261; 
@(negedge clk)
!rst && Lreq   ##1 !Lreq && !Nreq  &&   !Sreq  &&   !rst  &&   Ereq|-> ##1(!nextstate[0]);
endproperty

property property_n264; 
@(negedge clk)
!Wreq && !Sreq  &&   !rst  &&   Nreq   ##1 !Nreq && !Ereq  &&   !Wreq  &&   !Sreq  &&   !rst  &&   Lreq|-> ##1(!nextstate[0]);
endproperty

property property_n265; 
@(negedge clk)
!rst && Wreq   ##1 !Nreq && !Ereq  &&   !Wreq  &&   !Sreq  &&   !rst  &&   Lreq|-> ##1(!nextstate[0]);
endproperty


property property_n268; 
@(negedge clk)
!rst && Sreq   ##1 !Sreq && !rst  &&   Nreq |-> ##1(!nextstate[0]);
endproperty


property property_n279; 
@(negedge clk)
 Nreq  ##1 !Nreq && Lreq|-> ##1(nextstate[1]);
endproperty

property property_n281; 
@(negedge clk)
!Ereq && !Wreq   ##1 Nreq && Ereq|-> ##1(nextstate[1]);
endproperty


property property_n285; 
@(negedge clk)
!Lflit_id[0] && !Nflit_id[0]  &&   !Eflit_id[0]  &&   !Wflit_id[0]  &&   !Sflit_id[0]  &&   !Wreq  &&   !Sreq  &&   !rst   ##1 !Nflit_id[2] && !Eflit_id[2]  &&   !Wflit_id[2]  &&   !Sflit_id[2]  &&   !Ereq  &&   !Lflit_id[2]  &&   !rst  &&   Lreq  &&   Nreq |-> ##1(!nextstate[1]);
endproperty

property property_n287; 
@(negedge clk)
!Lreq && !Sreq  &&   !rst  &&   Lflit_id[0]   ##1 !Nflit_id[2] && !Eflit_id[2]  &&   !Wflit_id[2]  &&   !Sflit_id[2]  &&   !Lflit_id[2]  &&   !rst  &&   Lreq|-> ##1(!nextstate[1]);
endproperty

property property_n289; 
@(negedge clk)
 1  ##1 rst |-> ##1 (!nextstate[1]);
endproperty

property property_n290; 
@(negedge clk)
 rst  ##1 !rst |-> ##1 (!nextstate[1]);
endproperty

property property_n291; 
@(negedge clk)
!Lreq && !Wreq  &&   Nreq  &&   Ereq   ##1 !Lflit_id[1] |->  ##1 (nextstate[2]);
endproperty

property property_n292; 
@(negedge clk)
!Lreq && !Wreq  &&   Nreq   ##1 !Lflit_id[1]& Ereq|-> ##1(nextstate[2]);
endproperty

property property_n293; 
@(negedge clk)
!Lreq && !Wreq  &&   Nreq  &&   Ereq   ##1 !Nflit_id[1] |->  ##1 (nextstate[2]);
endproperty

property property_n294; 
@(negedge clk)
!Lreq && !Wreq  &&   Nreq   ##1 !Nflit_id[1]& Ereq|-> ##1(nextstate[2]);
endproperty

property property_n295; 
@(negedge clk)
!Lreq && !Wreq  &&   Nreq  &&   Ereq   ##1 !Eflit_id[1]|-> ##1 (nextstate[2]);
endproperty

property property_n296; 
@(negedge clk)
!Lreq && !Wreq  &&   Nreq   ##1 !Eflit_id[1]& Ereq|-> ##1(nextstate[2]);
endproperty

property property_n297; 
@(negedge clk)
!Lreq && !Wreq  &&   Nreq  &&   Ereq   ##1 !Wflit_id[1] |-> ##1 (nextstate[2]);
endproperty

property property_n298; 
@(negedge clk)
!Lreq && !Wreq  &&   Nreq   ##1 !Wflit_id[1] && Ereq |-> ##1(nextstate[2]);
endproperty

property property_n299; 
@(negedge clk)
!Lreq && !Wreq  &&   Nreq  &&   Ereq   ##1 !Sflit_id[1] |-> ##1 (nextstate[2]);
endproperty

property property_n300; 
@(negedge clk)
!Lreq && !Wreq  &&   Nreq   ##1 !Sflit_id[1] && Ereq |-> ##1(nextstate[2]);
endproperty

property property_n305; 
@(negedge clk)
 Lreq  ##1 !Lreq && Nreq |-> ##1(nextstate[2]);
endproperty

property property_n311; 
@(negedge clk)
!Ereq && !rst  &&   Lreq  &&   Nreq  &&   Wreq   ##1 !Nflit_id[2] && !Eflit_id[2]  &&   !Wflit_id[2]  &&   !Sflit_id[2]  &&   !Sreq  &&   !Lflit_id[2]  &&   !rst  &&   Lreq  &&   Nreq  &&   Ereq  &&   Wreq|-> ##1(!nextstate[2]);
endproperty

property property_n312; 
@(negedge clk)
!Sreq && !rst  &&   Lflit_id[0]  &&   Lreq  &&   Nreq  &&   Ereq  &&   Wreq   ##1 !Nflit_id[2] && !Eflit_id[2]  &&   !Wflit_id[2]  &&   !Sflit_id[2]  &&   !Sreq  &&   !Lflit_id[2]  &&   !rst  &&   Lreq  &&   Nreq  &&   Ereq  &&   Wreq|-> ##1(!nextstate[2]);
endproperty

property property_n313; 
@(negedge clk)
!Nreq && !rst   ##1 !rst && Lreq  &&   Nreq |-> ##1(!nextstate[2]);
endproperty

property property_n316; 
@(negedge clk)
 1  ##1 rst |-> ##1 (!nextstate[2]);
endproperty

property property_n317; 
@(negedge clk)
 rst  ##1 !rst |-> ##1 (!nextstate[2]);
endproperty

property property_n318; 
@(negedge clk)
!Lreq && Ereq   ##1 Lreq && Ereq|-> ##1(nextstate[3]);
endproperty


property property_n322; 
@(negedge clk)
!Lreq && !Sreq  &&   !rst  &&   Lflit_id[2]  &&   Nreq  &&   Ereq   ##1 !Nflit_id[2] && !Eflit_id[2]  &&   !Wflit_id[2]  &&   !Sflit_id[2]  &&   !Lreq  &&   !Sreq  &&   !Lflit_id[2]  &&   !rst  &&   Nreq  &&   Ereq|-> ##1(!nextstate[3]);
endproperty

property property_n323; 
@(negedge clk)
!Lreq && !Sreq  &&   !rst  &&   Nreq  &&   Ereq   ##1 !Lreq && !Sreq  &&   !rst  &&   Lflit_id[2]  &&   Nreq  &&   Ereq|-> ##1(!nextstate[3]);
endproperty

property property_n324; 
@(negedge clk)
!Nreq && !rst  &&   Lreq  &&   Ereq   ##1 !rst && Lreq  &&   Nreq  &&   Ereq|-> ##1(!nextstate[3]);
endproperty

property property_n325; 
@(negedge clk)
!Ereq && !rst   ##1 !rst && Nreq  &&   Ereq|-> ##1(!nextstate[3]);
endproperty

property property_n327; 
@(negedge clk)
 1  ##1 rst |-> ##1 (!nextstate[3]);
endproperty

property property_n328; 
@(negedge clk)
 rst  ##1 !rst |-> ##1 (!nextstate[3]);
endproperty

property property_n342; 
@(negedge clk)
 Ereq  ##1  !Ereq && Wreq|-> ##1(nextstate[4]);
endproperty

property property_n344; 
@(negedge clk)
!Ereq && !Wreq  &&   !rst  &&   Lflit_id[2]   ##1 !Ereq && !rst  &&   Wreq|-> ##1(!nextstate[4]);
endproperty

property property_n345; 
@(negedge clk)
!Wreq && !rst   ##1 !rst && Ereq  &&   Wreq|-> ##1(!nextstate[4]);
endproperty


property property_n347; 
@(negedge clk)
 1  ##1 rst |-> ##1 (!nextstate[4]);
endproperty

property property_n348; 
@(negedge clk)
 rst  ##1 !rst |-> ##1 (!nextstate[4]);
endproperty


property property_n350; 
@(negedge clk)
!Lflit_id[2] && !Nreq   ##1 !Nflit_id[1]& Nreq|-> ##2 (nextstate[0]);
endproperty

property property_n351; 
@(negedge clk)
!Lflit_id[2] && !Nreq   ##1 !Eflit_id[1]& Nreq|-> ##2 (nextstate[0]);
endproperty

property property_n352; 
@(negedge clk)
!Lflit_id[2] && !Nreq   ##1 !Wflit_id[1]& Nreq|-> ##2 (nextstate[0]);
endproperty

property property_n354; 
@(negedge clk)
!Lflit_id[1]& Sreq   ##1 !Sreq |-> ##1 ##1 (nextstate[0]);
endproperty


property property_n357; 
@(negedge clk)
!Lreq && !Nreq  &&   !Ereq  &&   !Wreq  &&   Lflit_id[2]   ##1 !Sreq |-> ##2  (nextstate[0]);
endproperty

property property_n358; 
@(negedge clk)
!Lreq && !Nreq  &&   !Ereq  &&   !Sreq  &&   Lflit_id[2]   ##1 !Wreq |-> ##2  (nextstate[0]);
endproperty

property property_n359; 
@(negedge clk)
!Lreq && !Nreq  &&   !Ereq  &&   Lflit_id[2]   ##1 !Wreq && !Sreq|-> ##2 (nextstate[0]);
endproperty

property property_n360; 
@(negedge clk)
!Lreq && !Nreq  &&   !Wreq  &&   !Sreq  &&   Lflit_id[2]   ##1 !Ereq |-> ##2  (nextstate[0]);
endproperty

property property_n361; 
@(negedge clk)
!Lreq && !Nreq  &&   !Wreq  &&   Lflit_id[2]   ##1  !Ereq && !Sreq|-> ##2 (nextstate[0]);
endproperty

property property_n362; 
@(negedge clk)
!Lreq && !Nreq  &&   !Sreq  &&   Lflit_id[2]   ##1 !Ereq && !Wreq|-> ##2 (nextstate[0]);
endproperty

property property_n363; 
@(negedge clk)
!Lreq && !Nreq  &&   Lflit_id[2]   ##1 !Ereq && !Wreq  &&   !Sreq|-> ##2 (nextstate[0]);
endproperty


property property_n366; 
@(negedge clk)
!Nreq && !Ereq  &&   !Wreq  &&   !Sreq  &&   Lflit_id[2]   ##1 !Lreq |-> ##2  (nextstate[0]);
endproperty

property property_n367; 
@(negedge clk)
!Nreq && !Ereq  &&   !Wreq  &&   Lflit_id[2]   ##1 !Lreq && !Sreq|-> ##2 (nextstate[0]);
endproperty

property property_n369; 
@(negedge clk)
!Nreq && !Ereq  &&   !Sreq  &&   Lflit_id[2]   ##1 !Lreq && !Wreq|-> ##2 (nextstate[0]);
endproperty

property property_n370; 
@(negedge clk)
!Nreq && !Ereq  &&   Lflit_id[2]   ##1 !Lreq && !Wreq  &&   !Sreq|-> ##2 (nextstate[0]);
endproperty

property property_n371; 
@(negedge clk)
!Nreq && !Wreq  &&   !Sreq  &&   Lflit_id[2]   ##1 !Lreq && !Ereq|-> ##2 (nextstate[0]);
endproperty

property property_n372; 
@(negedge clk)
!Nreq && !Wreq  &&   Lflit_id[2]   ##1 !Lreq && !Ereq  &&   !Sreq|-> ##2 (nextstate[0]);
endproperty

property property_n373; 
@(negedge clk)
!Nreq && !Sreq  &&   Lflit_id[2]   ##1 !Lreq && !Ereq  &&   !Wreq|-> ##2 (nextstate[0]);
endproperty

property property_n374; 
@(negedge clk)
!Nreq && Lflit_id[2]   ##1 !Lreq && !Ereq  &&   !Wreq  &&   !Sreq|-> ##2 (nextstate[0]);
endproperty

property property_n377; 
@(negedge clk)
!Sreq  ##1 !Lreq && Sreq|-> ##2 (nextstate[0]);
endproperty

property property_n378; 
@(negedge clk)
!Wreq && !Sreq  &&   Lreq  &&   Nreq   ##1 !Nreq |-> ##2  (nextstate[0]);
endproperty

property property_n379; 
@(negedge clk)
 1  ##1 rst |-> ##2  (nextstate[0]);
endproperty


property property_n381; 
@(negedge clk)
!Lflit_id[2] && !Lflit_id[1] &&   !Nflit_id[1] &&   !Eflit_id[1] &&   !Sflit_id[1] &&   !Wflit_id[1] &&   !rst  &&   Sreq   ##1 !Nflit_id[2] && !Eflit_id[2]  &&   !Wflit_id[2]  &&   !Sflit_id[2]  &&   !Lflit_id[2]  &&   !rst  &&   Sreq|-> ##2 (!nextstate[0]);
endproperty

property property_n382; 
@(negedge clk)
!Lreq && !Nreq  &&   !Sreq  &&   !rst  &&   Ereq  &&   Wreq   ##1 !Nflit_id[2] && !Eflit_id[2]  &&   !Wflit_id[2]  &&   !Sflit_id[2]  &&   !Lreq  &&   !Nreq  &&   !Sreq  &&   !Lflit_id[2]  &&   !rst  &&   Wreq|-> ##2 (!nextstate[0]);
endproperty

property property_n383; 
@(negedge clk)
!rst && Lflit_id[1] &&   Sreq   ##1 !Nflit_id[2] && !Eflit_id[2]  &&   !Wflit_id[2]  &&   !Sflit_id[2]  &&   !Lflit_id[2]  &&   !rst|-> ##2 (!nextstate[0]);
endproperty


property property_n385; 
@(negedge clk)
!Lreq && !Nreq  &&   !Wreq  &&   !Sreq  &&   !rst  &&   Lflit_id[2]  &&   Ereq   ##1 !Lreq && !Nreq  &&   !Wreq  &&   !Sreq  &&   !rst  &&   Ereq|-> ##2 (!nextstate[0]);
endproperty


property property_n387; 
@(negedge clk)
!Lreq && !Nreq  &&   !Sreq  &&   !rst  &&   Wreq   ##1 !Lreq && !Sreq  &&   !rst  &&   Nreq  &&   Wreq|-> ##2 (!nextstate[0]);
endproperty

property property_n388; 
@(negedge clk)
!Lreq && !Sreq  &&   !rst  &&   Nreq  &&   Wreq   ##1 !Lreq && !Sreq  &&   !rst  &&   Wreq|-> ##2 (!nextstate[0]);
endproperty

property property_n389; 
@(negedge clk)
!Lreq && !Wreq  &&   !Sreq  &&   !rst  &&   Nreq   ##1 !Nreq && !rst|-> ##2 (!nextstate[0]);
endproperty


property property_n391; 
@(negedge clk)
!Sreq && !rst  &&   Lreq  &&   Wreq   ##1 !Lreq && !Sreq  &&   !rst  &&   Wreq|-> ##2 (!nextstate[0]);
endproperty


property property_n393; 
@(negedge clk)
!Nreq && !Ereq  &&   !Wreq  &&   !Sreq  &&   !rst  &&   Lreq   ##1 !Nreq && !Ereq  &&   !Wreq  &&   !rst  &&   Lreq  &&   Sreq|-> ##2 (!nextstate[0]);
endproperty

property property_n394; 
@(negedge clk)
!Nreq && !Ereq  &&   !Wreq  &&   !Sreq  &&   !rst  &&   Lreq   ##1 !Nreq && !rst  &&   Lreq  &&   Ereq|-> ##2 (!nextstate[0]);
endproperty

property property_n395; 
@(negedge clk)
!Wreq && !Sreq  &&   !rst  &&   Lflit_id[0]   ##1 !Wreq && !Sreq  &&   !rst  &&   Nreq|-> ##2 (!nextstate[0]);
endproperty

property property_n396; 
@(negedge clk)
!Wreq && !Sreq  &&   !rst   ##1 !rst && Nreq  &&   Wreq|-> ##2 (!nextstate[0]);
endproperty

property property_n398; 
@(negedge clk)
!Sreq && !rst  &&   Wreq   ##1 !Sreq && !rst  &&   Lreq  &&   Wreq|-> ##2 (!nextstate[0]);
endproperty

property property_n399; 
@(negedge clk)
!Sreq && !rst  &&   Wreq   ##1 !rst && Sreq|-> ##2 (!nextstate[0]);
endproperty

property property_n401; 
@(negedge clk)
!Lflit_id[1] && !Wreq  &&   Lreq   ##1 Ereq |-> ##1 ##1 (nextstate[1]);
endproperty

property property_n402; 
@(negedge clk)
!Lflit_id[1] && !Wreq  &&   Ereq   ##1 Lreq |-> ##2 (nextstate[1]);
endproperty

property property_n403; 
@(negedge clk)
!Lflit_id[1] && !Wreq   ##1 Lreq && Ereq|-> ##2 (nextstate[1]);
endproperty

property property_n404; 
@(negedge clk)
!Lflit_id[1] && !Wreq  &&   Ereq  &&   Sreq   ##1 1 |-> ##2 (nextstate[1]);
endproperty

property property_n405; 
@(negedge clk)
!Lflit_id[1] && !Wreq  &&   Ereq   ##1 Sreq |-> ##2 (nextstate[1]);
endproperty

property property_n406; 
@(negedge clk)
!Lflit_id[1] && !Wreq  &&   Sreq   ##1 Ereq |-> ##2 (nextstate[1]);
endproperty

property property_n407; 
@(negedge clk)
!Lflit_id[1] && !Wreq   ##1 Ereq && Sreq|-> ##2 (nextstate[1]);
endproperty

property property_n408; 
@(negedge clk)
!Lreq  ##1 Ereq && Sreq|-> ##2 (nextstate[1]);
endproperty

property property_n409; 
@(negedge clk)
!Sreq && Lreq   ##1 !Ereq && Sreq|-> ##2 (nextstate[1]);
endproperty

property property_n410; 
@(negedge clk)
 Sreq  ##1 !Sreq && Lreq|-> ##2 (nextstate[1]);
endproperty

property property_n411; 
@(negedge clk)
!Lflit_id[2] && !Nflit_id[2]  &&   !Eflit_id[2]  &&   !Wflit_id[2]  &&   !Sflit_id[2]  &&   !Lreq  &&   !Nreq  &&   !Wreq  &&   !Sreq  &&   !rst  &&   Ereq   ##1 !Lflit_id[0] && !Nflit_id[0]  &&   !Eflit_id[0]  &&   !Wflit_id[0]  &&   !Sflit_id[0]  &&   !Lreq  &&   !Nreq  &&   !Wreq  &&   !Sreq  &&   !rst|-> ##2 (!nextstate[1]);
endproperty

property property_n412; 
@(negedge clk)
!Lflit_id[2] && !Nflit_id[2]  &&   !Eflit_id[2]  &&   !Wflit_id[2]  &&   !Sflit_id[2]  &&   !Lreq  &&   !Nreq  &&   !Wreq  &&   !Sreq  &&   !rst   ##1 !Lflit_id[0] && !Nflit_id[0]  &&   !Eflit_id[0]  &&   !Wflit_id[0]  &&   !Sflit_id[0]  &&   !Lreq  &&   !Wreq  &&   !Sreq  &&   !rst  &&   Nreq|-> ##2 (!nextstate[1]);
endproperty

property property_n413; 
@(negedge clk)
!Lflit_id[2] && !Nflit_id[2]  &&   !Eflit_id[2]  &&   !Wflit_id[2]  &&   !Sflit_id[2]  &&   !Lreq  &&   !Wreq  &&   !Sreq  &&   !rst  &&   Nreq   ##1 !Lflit_id[0] && !Nflit_id[0]  &&   !Eflit_id[0]  &&   !Wflit_id[0]  &&   !Sflit_id[0]  &&   !Lreq  &&   !Wreq  &&   !Sreq  &&   !rst  &&   Lflit_id[2]  &&   Nreq|-> ##2 (!nextstate[1]);
endproperty

property property_n414; 
@(negedge clk)
!Lflit_id[2] && !Nflit_id[2]  &&   !Eflit_id[2]  &&   !Wflit_id[2]  &&   !Sflit_id[2]  &&   !Lreq  &&   !Sreq  &&   !rst  &&   Wreq   ##1 !Lflit_id[0] && !Nflit_id[0]  &&   !Eflit_id[0]  &&   !Wflit_id[0]  &&   !Sflit_id[0]  &&   !Lreq  &&   !Wreq  &&   !Sreq  &&   !rst|-> ##2 (!nextstate[1]);
endproperty

property property_n415; 
@(negedge clk)
!Lflit_id[2] && !Nflit_id[2]  &&   !Eflit_id[2]  &&   !Wflit_id[2]  &&   !Sflit_id[2]  &&   !Lreq  &&   !Sreq  &&   !rst   ##1 !Lflit_id[0] && !Nflit_id[0]  &&   !Eflit_id[0]  &&   !Wflit_id[0]  &&   !Sflit_id[0]  &&   !Lreq  &&   !Sreq  &&   !rst  &&   Wreq|-> ##2 (!nextstate[1]);
endproperty

property property_n416; 
@(negedge clk)
!Lreq && !Ereq  &&   !rst   ##1 !Nflit_id[2] && !Eflit_id[2]  &&   !Wflit_id[2]  &&   !Sflit_id[2]  &&   !Ereq  &&   !Lflit_id[2]  &&   !rst  &&   Lreq  &&   Sreq|-> ##2 (!nextstate[1]);
endproperty

property property_n417; 
@(negedge clk)
!Nreq && !rst  &&   Lreq  &&   Ereq  &&   Sreq   ##1  !Nflit_id[2] && !Eflit_id[2]  &&   !Wflit_id[2]  &&   !Sflit_id[2]  &&   !Lflit_id[2]  &&   !rst  &&   Lreq  &&   Nreq  &&   Ereq  &&   Sreq|-> ##2 (!nextstate[1]);
endproperty

property property_n418; 
@(negedge clk)
!rst && Lreq  &&   Ereq  &&   Sreq   ##1 !Nflit_id[2] && !Eflit_id[2]  &&   !Wflit_id[2]  &&   !Sflit_id[2]  &&   !Nreq  &&   !Lflit_id[2]  &&   !rst  &&   Lreq  &&   Ereq  &&   Sreq|-> ##2 (!nextstate[1]);
endproperty

property property_n419; 
@(negedge clk)
!Ereq && !rst  &&   Lflit_id[2]  &&   Lreq  &&   Sreq   ##1 !Nflit_id[2] && !Eflit_id[2]  &&   !Wflit_id[2]  &&   !Sflit_id[2]  &&   !Ereq  &&   !Lflit_id[2]  &&   !rst  &&   Lreq  &&   Sreq|-> ##2 (!nextstate[1]);
endproperty

property property_n420; 
@(negedge clk)
!Ereq && !rst  &&   Lreq   ##1 !Nflit_id[2] && !Eflit_id[2]  &&   !Wflit_id[2]  &&   !Sflit_id[2]  &&   !Lflit_id[2]  &&   !rst  &&   Lreq  &&   Ereq  &&   Sreq|-> ##2 (!nextstate[1]);
endproperty

property property_n421; 
@(negedge clk)
!rst && Ereq   ##1 !Nflit_id[2] && !Eflit_id[2]  &&   !Wflit_id[2]  &&   !Sflit_id[2]  &&   !Ereq  &&   !Lflit_id[2]  &&   !rst  &&   Lreq  &&   Sreq|-> ##2 (!nextstate[1]);
endproperty

property property_n422; 
@(negedge clk)
!Lreq && !Sreq  &&   !rst  &&   Lflit_id[2]   ##1 !Lreq && !Sreq  &&   !rst|-> ##2 (!nextstate[1]);
endproperty

property property_n423; 
@(negedge clk)
!Lreq && !rst  &&   Sreq   ##1 !Lreq && !Sreq  &&   !rst|-> ##2 (!nextstate[1]);
endproperty

property property_n424; 
@(negedge clk)
!Lreq && !rst   ##1 !Lreq && !rst  &&   Sreq|-> ##2 (!nextstate[1]);
endproperty

property property_n425; 
@(negedge clk)
!rst && Lreq   ##1 !Lreq && !rst|-> ##2 (!nextstate[1]);
endproperty

property property_n428; 
@(negedge clk)
!Lreq && Nreq   ##1 Lreq && Wreq|-> ##2 (nextstate[2]);
endproperty

property property_n431; 
@(negedge clk)
 Lreq  ##1 !Lreq && Nreq|-> ##2 (nextstate[2]);
endproperty

property property_n432; 
@(negedge clk)
!Lflit_id[2] && !Lflit_id[1] &&   !Nflit_id[2]  &&   !Eflit_id[2]  &&   !Wflit_id[2]  &&   !Sflit_id[2]  &&   !Wreq  &&   !rst  &&   Lreq  &&   Nreq   ##1 !Lflit_id[0] && !Nflit_id[0]  &&   !Eflit_id[0]  &&   !Wflit_id[0]  &&   !Sflit_id[0]  &&   !Wreq  &&   !rst  &&   Lreq  &&   Nreq|-> ##2 (!nextstate[2]);
endproperty

property property_n435; 
@(negedge clk)
!Lflit_id[2] && !Nflit_id[2]  &&   !Eflit_id[2]  &&   !Wflit_id[2]  &&   !Sflit_id[2]  &&   !Nreq  &&   !Sreq  &&   !rst   ##1 !Lflit_id[0] && !Nflit_id[0]  &&   !Eflit_id[0]  &&   !Wflit_id[0]  &&   !Sflit_id[0]  &&   !Nreq  &&   !rst  &&   Sreq|-> ##2 (!nextstate[2]);
endproperty

property property_n436; 
@(negedge clk)
!Lflit_id[2] && !Nflit_id[2]  &&   !Eflit_id[2]  &&   !Wflit_id[2]  &&   !Sflit_id[2]  &&   !Nreq  &&   !rst  &&   Sreq   ##1 !Lflit_id[0] && !Nflit_id[0]  &&   !Eflit_id[0]  &&   !Wflit_id[0]  &&   !Sflit_id[0]  &&   !Nreq  &&   !rst|-> ##2 (!nextstate[2]);
endproperty

property property_n437; 
@(negedge clk)
!Lflit_id[2] && !Nflit_id[2]  &&   !Eflit_id[2]  &&   !Wflit_id[2]  &&   !Sflit_id[2]  &&   !Ereq  &&   !rst  &&   Lreq  &&   Nreq  &&   Wreq  &&   Sreq   ##1 !Lflit_id[0] && !Nflit_id[0]  &&   !Eflit_id[0]  &&   !Wflit_id[0]  &&   !Sflit_id[0]  &&   !rst  &&   Lflit_id[2]  &&   Lreq  &&   Nreq  &&   Wreq|-> ##2 (!nextstate[2]);
endproperty

property property_n438; 
@(negedge clk)
!Lflit_id[2] && !Lreq  &&   !Nreq  &&   !Sreq  &&   !rst   ##1 !Lreq && !Sreq  &&   !rst  &&   Nreq|-> ##2 (!nextstate[2]);
endproperty

property property_n439; 
@(negedge clk)
!Lreq && !rst  &&   Nreq   ##1 !Wreq && !rst  &&   Lreq  &&   Nreq|-> ##2 (!nextstate[2]);
endproperty

property property_n440; 
@(negedge clk)
!Nreq && !rst  &&   Lflit_id[2]   ##1 !Nreq && !rst|-> ##2 (!nextstate[2]);
endproperty

property property_n441; 
@(negedge clk)
!Nreq && !rst   ##1 !rst && Lreq  &&   Nreq|-> ##2 (!nextstate[2]);
endproperty

property property_n442; 
@(negedge clk)
!rst && Nreq   ##1 !Nreq && !rst|-> ##2 (!nextstate[2]);
endproperty

property property_n443; 
@(negedge clk)
!Wreq && !rst  &&   Lflit_id[2]  &&   Lreq  &&   Nreq   ##1 !Wreq && !rst  &&   Lreq  &&   Nreq|-> ##2 (!nextstate[2]);
endproperty

property property_n444; 
@(negedge clk)
 1  ##1 rst |-> ##2 (!nextstate[2]);
endproperty

property property_n445; 
@(negedge clk)
 rst  ##1 !rst |-> ##2 (!nextstate[2]);
endproperty

property property_n446; 
@(negedge clk)
!Lreq && Ereq   ##1  Lreq && Ereq|-> ##2 (nextstate[3]);
endproperty

property property_n447; 
@(negedge clk)
!Nreq && !Wreq  &&   Lreq   ##1 Ereq |-> ##2 (nextstate[3]);
endproperty

property property_n448; 
@(negedge clk)
!Nreq && !Sreq  &&   Lreq   ##1 Ereq |-> ##2 (nextstate[3]);
endproperty

property property_n449; 
@(negedge clk)
!Wreq && Lflit_id[2]   ##1 !Nreq && Ereq|-> ##2 (nextstate[3]);
endproperty

property property_n450; 
@(negedge clk)
!Wreq && Lreq   ##1 !Nreq && Ereq|-> ##2 (nextstate[3]);
endproperty

property property_n451; 
@(negedge clk)
 Lflit_id[2]  ##1 !Nreq && !Wreq  &&   Ereq|-> ##2 (nextstate[3]);
endproperty


property property_n453; 
@(negedge clk)
!Sreq && Lreq   ##1 !Nreq && Ereq|-> ##2 (nextstate[3]);
endproperty

property property_n454; 
@(negedge clk)
 Nreq  ##1 !Nreq && Ereq|-> ##2 (nextstate[3]);
endproperty

property property_n455; 
@(negedge clk)
!Lflit_id[2] && !Nflit_id[2]  &&   !Eflit_id[2]  &&   !Wflit_id[2]  &&   !Sflit_id[2]  &&   !Lreq  &&   !Sreq  &&   !rst  &&   Nreq  &&   Ereq   ##1 !Lflit_id[0] && !Nflit_id[0]  &&   !Eflit_id[0]  &&   !Wflit_id[0]  &&   !Sflit_id[0]  &&   !Lreq  &&   !Sreq  &&   !rst  &&   Lflit_id[2]  &&   Nreq  &&   Ereq|-> ##2 (!nextstate[3]);
endproperty

property property_n456; 
@(negedge clk)
!Lflit_id[0] && !Nflit_id[0]  &&   !Eflit_id[0]  &&   !Wflit_id[0]  &&   !Sflit_id[0]  &&   !Wreq  &&   !rst  &&   Lreq  &&   Nreq  &&   Ereq  &&   Sreq   ##1  !Lflit_id[1]& !Nflit_id[1] &&   !Eflit_id[1] &&   !Wflit_id[1] &&   !Sflit_id[1] &&   !rst  &&   Lreq  &&   Nreq  &&   Ereq  &&   Sreq|-> ##2 (!nextstate[3]);
endproperty

property property_n457; 
@(negedge clk)
!Lflit_id[0] && !Nflit_id[0]  &&   !Eflit_id[0]  &&   !Wflit_id[0]  &&   !Sflit_id[0]  &&   !Sreq  &&   !rst  &&   Lflit_id[2]  &&   Lreq  &&   Nreq  &&   Ereq   ##1  !Lflit_id[1]& !Nflit_id[1] &&   !Eflit_id[1] &&   !Wflit_id[1] &&   !Sflit_id[1] &&   !Sreq  &&   !rst  &&   Lreq  &&   Nreq  &&   Ereq|-> ##2 (!nextstate[3]);
endproperty

property property_n458; 
@(negedge clk)
!Lflit_id[0] && !Nflit_id[0]  &&   !Eflit_id[0]  &&   !Wflit_id[0]  &&   !Sflit_id[0]  &&   !Lreq  &&   !Nreq  &&   !Ereq  &&   !Wreq  &&   !Sreq  &&   !rst   ##1  !Nflit_id[2] && !Eflit_id[2]  &&   !Wflit_id[2]  &&   !Sflit_id[2]  &&   !Lreq  &&   !Ereq  &&   !Wreq  &&   !Sreq  &&   !Lflit_id[2]  &&   !rst|-> ##2 (!nextstate[3]);
endproperty

property property_n459; 
@(negedge clk)
!Lflit_id[0] && !Nflit_id[0]  &&   !Eflit_id[0]  &&   !Wflit_id[0]  &&   !Sflit_id[0]  &&   !Lreq  &&   !Ereq  &&   !Wreq  &&   !Sreq  &&   !rst   ##1 !Nflit_id[2] && !Eflit_id[2]  &&   !Wflit_id[2]  &&   !Sflit_id[2]  &&   !Lreq  &&   !Ereq  &&   !Wreq  &&   !Lflit_id[2]  &&   !rst  &&   Sreq|-> ##2 (!nextstate[3]);
endproperty

property property_n460; 
@(negedge clk)
!Lflit_id[0] && !Nflit_id[0]  &&   !Eflit_id[0]  &&   !Wflit_id[0]  &&   !Sflit_id[0]  &&   !Lreq  &&   !Ereq  &&   !Wreq  &&   !rst  &&   Sreq   ##1 !Nflit_id[2] && !Eflit_id[2]  &&   !Wflit_id[2]  &&   !Sflit_id[2]  &&   !Lreq  &&   !Ereq  &&   !Wreq  &&   !Lflit_id[2]  &&   !rst|-> ##2 (!nextstate[3]);
endproperty

property property_n461; 
@(negedge clk)
!Lflit_id[0] && !Nflit_id[0]  &&   !Eflit_id[0]  &&   !Wflit_id[0]  &&   !Sflit_id[0]  &&   !Lreq  &&   !Ereq  &&   !Wreq  &&   !rst   ##1 !Nflit_id[2] && !Eflit_id[2]  &&   !Wflit_id[2]  &&   !Sflit_id[2]  &&   !Ereq  &&   !Wreq  &&   !Lflit_id[2]  &&   !rst  &&   Lreq|-> ##2 (!nextstate[3]);
endproperty

property property_n462; 
@(negedge clk)
!Lflit_id[0] && !Nflit_id[0]  &&   !Eflit_id[0]  &&   !Wflit_id[0]  &&   !Sflit_id[0]  &&   !Ereq  &&   !Wreq  &&   !rst  &&   Lreq   ##1 !Nflit_id[2] && !Eflit_id[2]  &&   !Wflit_id[2]  &&   !Sflit_id[2]  &&   !Lreq  &&   !Ereq  &&   !Wreq  &&   !Lflit_id[2]  &&   !rst|-> ##2 (!nextstate[3]);
endproperty

property property_n463; 
@(negedge clk)
!Lflit_id[0] && !Nflit_id[0]  &&   !Eflit_id[0]  &&   !Wflit_id[0]  &&   !Sflit_id[0]  &&   !Ereq  &&   !Wreq  &&   !rst  &&   Lflit_id[2]  &&   Lreq   ##1 !Nflit_id[2] && !Eflit_id[2]  &&   !Wflit_id[2]  &&   !Sflit_id[2]  &&   !Ereq  &&   !Wreq  &&   !Lflit_id[2]  &&   !rst  &&   Lreq|-> ##2 (!nextstate[3]);
endproperty

property property_n464; 
@(negedge clk)
!Ereq && !Wreq  &&   !rst  &&   Lflit_id[0]   ##1 !Nflit_id[2] && !Eflit_id[2]  &&   !Wflit_id[2]  &&   !Sflit_id[2]  &&   !Ereq  &&   !Wreq  &&   !Lflit_id[2]  &&   !rst|-> ##2 (!nextstate[3]);
endproperty

property property_n465; 
@(negedge clk)
!Ereq && !Wreq  &&   !rst   ##1 !Nflit_id[2] && !Eflit_id[2]  &&   !Wflit_id[2]  &&   !Sflit_id[2]  &&   !Ereq  &&   !Lflit_id[2]  &&   !rst  &&   Wreq |-> ##2 (!nextstate[3]);
endproperty

property property_n466; 
@(negedge clk)
!Ereq && !rst  &&   Wreq   ##1 !Nflit_id[2] && !Eflit_id[2]  &&   !Wflit_id[2]  &&   !Sflit_id[2]  &&   !Ereq  &&   !Lflit_id[2]  &&   !rst |-> ##2 (!nextstate[3]);
endproperty

property property_n467; 
@(negedge clk)
!Lreq && !Nreq  &&   !Sreq  &&   !rst  &&   Ereq   ##1 !Lreq && !Sreq  &&   !rst  &&   Nreq  &&   Ereq|-> ##2 (!nextstate[3]);
endproperty


property property_n469; 
@(negedge clk)
!Lreq && !Nreq  &&   !Ereq  &&   !Wreq  &&   !Sreq  &&   !rst   ##1 !Nreq && !rst  &&   Ereq|-> ##2 (!nextstate[3]);
endproperty

property property_n470; 
@(negedge clk)
!Nreq && !Ereq  &&   !rst  &&   Wreq   ##1 !Nreq && !rst  &&   Ereq|-> ##2 (!nextstate[3]);
endproperty

property property_n471; 
@(negedge clk)
!Nreq && !rst  &&   Lreq  &&   Ereq   ##1 !rst && Lreq  &&   Nreq  &&   Ereq|-> ##2 (!nextstate[3]);
endproperty



property property_n473; 
@(negedge clk)
!Ereq && !rst   ##1 !rst && Nreq  &&   Ereq|-> ##2 (!nextstate[3]);
endproperty

property property_n474; 
@(negedge clk)
!rst && Ereq   ##1 !Ereq && !rst|-> ##2 (!nextstate[3]);
endproperty

property property_n475; 
@(negedge clk)
 1  ##1 rst |-> ##2 (!nextstate[3]);
endproperty

property property_n476; 
@(negedge clk)
rst  ##1 !rst |-> ##2 (!nextstate[3]);
endproperty

property property_n477; 
@(negedge clk)
!Ereq && Wreq   ##1 !Lflit_id[1]& Ereq|-> ##2 (nextstate[4]);
endproperty

property property_n478; 
@(negedge clk)
!Ereq && Lflit_id[2]  &&   Sreq   ##1 Wreq |-> ##2 (nextstate[4]);
endproperty

property property_n480; 
@(negedge clk)
Lflit_id[2] && Sreq   ##1 !Ereq && Wreq|-> ##2 (nextstate[4]);
endproperty


property property_n482; 
@(negedge clk)
Ereq  ##1 !Ereq && Wreq|-> ##2 (nextstate[4]);
endproperty

property property_n483; 
@(negedge clk)
!Lflit_id[2] && !Nflit_id[2]  &&   !Eflit_id[2]  &&   !Wflit_id[2]  &&   !Sflit_id[2]  &&   !Wreq  &&   !rst   ##1 !Lflit_id[0] && !Nflit_id[0]  &&   !Eflit_id[0]  &&   !Wflit_id[0]  &&   !Sflit_id[0]  &&   !Wreq  &&   !rst  &&   Lflit_id[2]|-> ##2 (!nextstate[4]);
endproperty

property property_n484; 
@(negedge clk)
!Ereq && !Wreq  &&   !Sreq  &&   !rst   ##1 !Nflit_id[2] && !Eflit_id[2]  &&   !Wflit_id[2]  &&   !Sflit_id[2]  &&   !Ereq  &&   !Lflit_id[2]  &&   !rst  &&   Wreq|-> ##2 (!nextstate[4]);
endproperty


property property_n486; 
@(negedge clk)
!Wreq && !rst   ##1 !rst && Ereq  &&   Wreq|-> ##2 (!nextstate[4]);
endproperty

property property_n487; 
@(negedge clk)
!rst && Wreq   ##1 !Wreq && !rst|-> ##2 (!nextstate[4]);
endproperty

property property_n488; 
@(negedge clk)
1  ##1 rst |-> ##2 (!nextstate[4]);
endproperty

property property_n489; 
@(negedge clk)
rst  ##1 !rst |-> ##2 (!nextstate[4]);
endproperty

property_0_assert : assert property (property_0) else $error("property_0 not held!");
property_1_assert : assert property (property_1) else $error("property_1 not held!");
property_2_assert : assert property (property_2) else $error("property_2  not held!");
property_3_assert : assert property (property_3) else $error("property_3 not held!");
property_4_assert : assert property (property_4) else $error("property_4 not held!");
property_5_assert : assert property (property_5) else $error("property_5 not held!");
property_6_assert : assert property (property_6) else $error("property_6 not held!");
property_7_assert : assert property (property_7) else $error("property_7 not held!");
property_8_assert : assert property (property_8) else $error("property_8 not held!");
property_9_assert : assert property (property_9) else $error("property_9 not held!");
property_10_assert : assert property (property_10) else $error("property_10 not held!");
property_11_assert : assert property (property_11) else $error("property_11 not held!");
property_12_assert : assert property (property_12) else $error("property_12 not held!");
property_13_assert : assert property (property_13) else $error("property_13 not held!");
property_14_assert : assert property (property_14) else $error("property_14 not held!");
property_15_assert : assert property (property_15) else $error("property_15 not held!");
property_16_assert : assert property (property_16) else $error("property_16 not held!");
property_17_assert : assert property (property_17) else $error("property_17 not held!");
property_18_assert : assert property (property_18) else $error("property_18 not held!");
property_19_assert : assert property (property_19) else $error("property_19 not held!");
property_20_assert : assert property (property_20) else $error("property_20 not held!");
property_21_assert : assert property (property_21) else $error("property_21 not held!");
property_22_assert : assert property (property_22) else $error("property_22 not held!");
property_23_assert : assert property (property_23) else $error("property_23 not held!");
property_24_assert : assert property (property_24) else $error("property_24 not held!");
property_25_assert : assert property (property_25) else $error("property_25 not held!");
property_26_assert : assert property (property_26) else $error("property_26 not held!");
property_27_assert : assert property (property_27) else $error("property_27 not held!");
property_28_assert : assert property (property_28) else $error("property_28 not held!");
property_29_assert : assert property (property_29) else $error("property_29 not held!");
property_30_assert : assert property (property_30) else $error("property_30 not held!");
property_31_assert : assert property (property_31) else $error("property_31 not held!");
property_32_assert : assert property (property_32) else $error("property_32 not held!");
property_33_assert : assert property (property_33) else $error("property_33 not held!");
property_34_assert : assert property (property_34) else $error("property_34 not held!");
property_35_assert : assert property (property_35) else $error("property_35 not held!");
property_36_assert : assert property (property_36) else $error("property_36 not held!");
property_37_assert : assert property (property_37) else $error("property_37 not held!");
property_38_assert : assert property (property_38) else $error("property_38 not held!");
property_39_assert : assert property (property_39) else $error("property_39 not held!");
property_40_assert : assert property (property_40) else $error("property_40 not held!");
property_41_assert : assert property (property_41) else $error("property_41 not held!");
property_42_assert : assert property (property_42) else $error("property_42 not held!");
property_43_assert : assert property (property_43) else $error("property_43 not held!");
property_44_assert : assert property (property_44) else $error("property_44 not held!");
property_45_assert : assert property (property_45) else $error("property_45 not held!");
property_46_assert : assert property (property_46) else $error("property_46 not held! ");
property_47_assert : assert property (property_47) else $error("property_47 not held! ");
property_48_assert : assert property (property_48) else $error("property_48 not held! ");
property_49_assert : assert property (property_49) else $error("property_49 not held! ");
property_50_assert : assert property (property_50) else $error("property_50 not held! ");
property_51_assert : assert property (property_51) else $error("property_51 not held! ");
property_52_assert : assert property (property_52) else $error("property_52 not held! ");
property_53_assert : assert property (property_53) else $error("property_53 not held! ");
property_54_assert : assert property (property_54) else $error("property_54 not held! ");
property_55_assert : assert property (property_55) else $error("property_55 not held! ");
property_56_assert : assert property (property_56) else $error("property_56 not held! ");
property_57_assert : assert property (property_57) else $error("property_57 not held! ");
property_58_assert : assert property (property_58) else $error("property_58 not held! ");
property_59_assert : assert property (property_59) else $error("property_59 not held! ");
property_60_assert : assert property (property_60) else $error("property_60 not held! ");
property_61_assert : assert property (property_61) else $error("property_61 not held! ");
property_62_assert : assert property (property_62) else $error("property_62 not held! ");
property_63_assert : assert property (property_63) else $error("property_63 not held! ");
property_64_assert : assert property (property_64) else $error("property_64 not held! ");
property_65_assert : assert property (property_65) else $error("property_65 not held! ");
property_66_assert : assert property (property_66) else $error("property_66 not held! ");
property_67_assert : assert property (property_67) else $error("property_67 not held! ");
property_68_assert : assert property (property_68) else $error("property_68 not held! ");
property_69_assert : assert property (property_69) else $error("property_69 not held! ");
property_70_assert : assert property (property_70) else $error("property_70 not held! ");
property_71_assert : assert property (property_71) else $error("property_71 not held! ");
property_72_assert : assert property (property_72) else $error("property_72 not held! ");
property_76_assert : assert property (property_76) else $error("property_76 not held! ");
property_77_assert : assert property (property_77) else $error("property_77 not held! ");
property_79_assert : assert property (property_79) else $error("property_79 not held! ");
property_80_assert : assert property (property_80) else $error("property_80 not held! ");
property_82_assert : assert property (property_82) else $error("property_82 not held! ");
property_83_assert : assert property (property_83) else $error("property_83 not held! ");
property_84_assert : assert property (property_84) else $error("property_84 not held! ");
property_86_assert : assert property (property_86) else $error("property_86 not held! ");
property_92_assert : assert property (property_92) else $error("property_92 not held! ");
property_93_assert : assert property (property_93) else $error("property_93 not held! ");
property_96_assert : assert property (property_96) else $error("property_96 not held! ");
property_98_assert : assert property (property_98) else $error("property_98 not held! ");
property_99_assert : assert property (property_99) else $error("property_99 not held! ");
property_100_assert : assert property (property_100) else $error("property_100 not held! ");
property_102_assert : assert property (property_102) else $error("property_102 not held! ");
property_103_assert : assert property (property_103) else $error("property_103 not held! ");
property_105_assert : assert property (property_105) else $error("property_105 not held! ");
property_106_assert : assert property (property_106) else $error("property_106 not held! ");
property_108_assert : assert property (property_108) else $error("property_108 not held! ");
property_109_assert : assert property (property_109) else $error("property_109 not held! ");
property_112_assert : assert property (property_112) else $error("property_112 not held! ");
property_114_assert : assert property (property_114) else $error("property_114 not held! ");
property_115_assert : assert property (property_115) else $error("property_115 not held! ");
property_117_assert : assert property (property_117) else $error("property_117 not held! ");
property_118_assert : assert property (property_118) else $error("property_118 not held! ");
property_121_assert : assert property (property_121) else $error("property_121 not held! ");
property_122_assert : assert property (property_122) else $error("property_122 not held! ");
property_123_assert : assert property (property_123) else $error("property_123 not held! ");
property_124_assert : assert property (property_124) else $error("property_124 not held! ");
property_125_assert : assert property (property_125) else $error("property_125 not held! ");
property_126_assert : assert property (property_126) else $error("property_126 not held! ");
property_127_assert : assert property (property_127) else $error("property_127 not held! ");
property_128_assert : assert property (property_128) else $error("property_128 not held! ");
property_129_assert : assert property (property_129) else $error("property_129 not held! ");
property_130_assert : assert property (property_130) else $error("property_130 not held! ");
property_131_assert : assert property (property_131) else $error("property_131 not held! ");
property_132_assert : assert property (property_132) else $error("property_132 not held! ");
property_133_assert : assert property (property_133) else $error("property_133 not held! ");
property_134_assert : assert property (property_134) else $error("property_134 not held! ");
property_135_assert : assert property (property_135) else $error("property_135 not held! ");
property_136_assert : assert property (property_136) else $error("property_136 not held! ");
property_137_assert : assert property (property_137) else $error("property_137 not held! ");
property_138_assert : assert property (property_138) else $error("property_138 not held! ");
property_139_assert : assert property (property_139) else $error("property_139 not held! ");
property_140_assert : assert property (property_140) else $error("property_140 not held! ");
property_141_assert : assert property (property_141) else $error("property_141 not held! ");
property_142_assert : assert property (property_142) else $error("property_142 not held! ");
property_143_assert : assert property (property_143) else $error("property_143 not held! ");
property_144_assert : assert property (property_144) else $error("property_144 not held! ");
property_145_assert : assert property (property_145) else $error("property_145 not held! ");
property_146_assert : assert property (property_146) else $error("property_146 not held! ");
property_147_assert : assert property (property_147) else $error("property_147 not held! ");
property_148_assert : assert property (property_148) else $error("property_148 not held! ");
property_149_assert : assert property (property_149) else $error("property_149 not held! ");
property_150_assert : assert property (property_150) else $error("property_150 not held! ");
property_152_assert : assert property (property_152) else $error("property_152 not held! ");
property_153_assert : assert property (property_153) else $error("property_153 not held! ");
property_154_assert : assert property (property_154) else $error("property_154 not held! ");
property_155_assert : assert property (property_155) else $error("property_155 not held! ");
property_156_assert : assert property (property_156) else $error("property_156 not held! ");
property_157_assert : assert property (property_157) else $error("property_157 not held! ");
property_158_assert : assert property (property_158) else $error("property_158 not held! ");
property_159_assert : assert property (property_159) else $error("property_159 not held! ");
property_160_assert : assert property (property_160) else $error("property_160 not held! ");
property_162_assert : assert property (property_162) else $error("property_162 not held! ");
property_163_assert : assert property (property_163) else $error("property_163 not held! ");
property_164_assert : assert property (property_164) else $error("property_164 not held! ");
property_165_assert : assert property (property_165) else $error("property_165 not held! ");
property_166_assert : assert property (property_166) else $error("property_166 not held! ");
property_167_assert : assert property (property_167) else $error("property_167 not held! ");
property_168_assert : assert property (property_168) else $error("property_168 not held! ");
property_169_assert : assert property (property_169) else $error("property_169 not held! ");
property_170_assert : assert property (property_170) else $error("property_170 not held! ");
property_171_assert : assert property (property_171) else $error("property_171 not held! ");
property_172_assert : assert property (property_172) else $error("property_172 not held! ");
property_173_assert : assert property (property_173) else $error("property_173 not held! ");
property_174_assert : assert property (property_174) else $error("property_174 not held! ");
property_175_assert : assert property (property_175) else $error("property_175 not held! ");
property_176_assert : assert property (property_176) else $error("property_176 not held! ");
property_177_assert : assert property (property_177) else $error("property_177 not held! ");
property_178_assert : assert property (property_178) else $error("property_178 not held! ");
property_179_assert : assert property (property_179) else $error("property_179 not held! ");
property_180_assert : assert property (property_180) else $error("property_180 not held! ");
property_181_assert : assert property (property_181) else $error("property_181 not held! ");
property_182_assert : assert property (property_182) else $error("property_182 not held! ");
property_183_assert : assert property (property_183) else $error("property_183 not held! ");
property_184_assert : assert property (property_184) else $error("property_184 not held! ");
property_185_assert : assert property (property_185) else $error("property_185 not held! ");
property_186_assert : assert property (property_186) else $error("property_186 not held! ");
property_187_assert : assert property (property_187) else $error("property_187 not held! ");
property_188_assert : assert property (property_188) else $error("property_188 not held! ");
property_190_assert : assert property (property_190) else $error("property_190 not held! ");

property_n1_assert : assert property (property_n1) else $error("property_n1 not held! ");
property_n2_assert : assert property (property_n2) else $error("property_n2 not held! ");
property_n3_assert : assert property (property_n3) else $error("property_n3 not held! ");
property_n4_assert : assert property (property_n4) else $error("property_n4 not held! ");
property_n5_assert : assert property (property_n5) else $error("property_n5 not held! ");
property_n6_assert : assert property (property_n6) else $error("property_n6 not held! ");
property_n7_assert : assert property (property_n7) else $error("property_n7 not held! ");
property_n8_assert : assert property (property_n8) else $error("property_n8 not held! ");
property_n9_assert : assert property (property_n9) else $error("property_n9 not held! ");
property_n10_assert : assert property (property_n10) else $error("property_n10 not held! ");
property_n11_assert : assert property (property_n11) else $error("property_n11 not held! ");
property_n12_assert : assert property (property_n12) else $error("property_n12 not held! ");
property_n13_assert : assert property (property_n13) else $error("property_n13 not held! ");
property_n14_assert : assert property (property_n14) else $error("property_n14 not held! ");
property_n15_assert : assert property (property_n15) else $error("property_n15 not held! ");
property_n16_assert : assert property (property_n16) else $error("property_n16 not held! ");
property_n17_assert : assert property (property_n17) else $error("property_n17 not held! ");
property_n18_assert : assert property (property_n18) else $error("property_n18 not held! ");
property_n19_assert : assert property (property_n19) else $error("property_n19 not held! ");
property_n20_assert : assert property (property_n20) else $error("property_n20 not held! ");
property_n21_assert : assert property (property_n21) else $error("property_n21 not held! ");
property_n22_assert : assert property (property_n22) else $error("property_n22 not held! ");
property_n23_assert : assert property (property_n23) else $error("property_n23 not held! ");
property_n24_assert : assert property (property_n24) else $error("property_n24 not held! ");
property_n25_assert : assert property (property_n25) else $error("property_n25 not held! ");
property_n26_assert : assert property (property_n26) else $error("property_n26 not held! ");
property_n27_assert : assert property (property_n27) else $error("property_n27 not held! ");
property_n28_assert : assert property (property_n28) else $error("property_n28 not held! ");
property_n29_assert : assert property (property_n29) else $error("property_n29 not held! ");
property_n30_assert : assert property (property_n30) else $error("property_n30 not held! ");
property_n31_assert : assert property (property_n31) else $error("property_n31 not held! ");
property_n32_assert : assert property (property_n32) else $error("property_n32 not held! ");
property_n33_assert : assert property (property_n33) else $error("property_n33 not held! ");
property_n34_assert : assert property (property_n34) else $error("property_n34 not held! ");
property_n35_assert : assert property (property_n35) else $error("property_n35 not held! ");
property_n36_assert : assert property (property_n36) else $error("property_n36 not held! ");
property_n37_assert : assert property (property_n37) else $error("property_n37 not held! ");
property_n38_assert : assert property (property_n38) else $error("property_n38 not held! ");
property_n39_assert : assert property (property_n39) else $error("property_n39 not held! ");
property_n40_assert : assert property (property_n40) else $error("property_n40 not held! ");
property_n41_assert : assert property (property_n41) else $error("property_n41 not held! ");
property_n42_assert : assert property (property_n42) else $error("property_n42 not held! ");
property_n43_assert : assert property (property_n43) else $error("property_n43 not held! ");
property_n44_assert : assert property (property_n44) else $error("property_n44 not held! ");
property_n45_assert : assert property (property_n45) else $error("property_n45 not held! ");
property_n46_assert : assert property (property_n46) else $error("property_n46 not held! ");
property_n47_assert : assert property (property_n47) else $error("property_n47 not held! ");
property_n48_assert : assert property (property_n48) else $error("property_n48 not held! ");
property_n49_assert : assert property (property_n49) else $error("property_n49 not held! ");
property_n50_assert : assert property (property_n50) else $error("property_n50 not held! ");
property_n51_assert : assert property (property_n51) else $error("property_n51 not held! ");
property_n52_assert : assert property (property_n52) else $error("property_n52 not held! ");
property_n53_assert : assert property (property_n53) else $error("property_n53 not held! ");
property_n54_assert : assert property (property_n54) else $error("property_n54 not held! ");
property_n55_assert : assert property (property_n55) else $error("property_n55 not held! ");
property_n56_assert : assert property (property_n56) else $error("property_n56 not held! ");
property_n57_assert : assert property (property_n57) else $error("property_n57 not held! ");
property_n58_assert : assert property (property_n58) else $error("property_n58 not held! ");
property_n59_assert : assert property (property_n59) else $error("property_n59 not held! ");
property_n60_assert : assert property (property_n60) else $error("property_n60 not held! ");
property_n61_assert : assert property (property_n61) else $error("property_n61 not held! ");
property_n62_assert : assert property (property_n62) else $error("property_n62 not held! ");
property_n63_assert : assert property (property_n63) else $error("property_n63 not held! ");
property_n64_assert : assert property (property_n64) else $error("property_n64 not held! ");
property_n65_assert : assert property (property_n65) else $error("property_n65 not held! ");
property_n66_assert : assert property (property_n66) else $error("property_n66 not held! ");
property_n67_assert : assert property (property_n67) else $error("property_n67 not held! ");
property_n68_assert : assert property (property_n68) else $error("property_n68 not held! ");
property_n69_assert : assert property (property_n69) else $error("property_n69 not held! ");
property_n70_assert : assert property (property_n70) else $error("property_n70 not held! ");
property_n71_assert : assert property (property_n71) else $error("property_n71 not held! ");
property_n72_assert : assert property (property_n72) else $error("property_n72 not held! ");
property_n73_assert : assert property (property_n73) else $error("property_n73 not held! ");
property_n74_assert : assert property (property_n74) else $error("property_n74 not held! ");
property_n75_assert : assert property (property_n75) else $error("property_n75 not held! ");
property_n76_assert : assert property (property_n76) else $error("property_n76 not held! ");
property_n77_assert : assert property (property_n77) else $error("property_n77 not held! ");
property_n78_assert : assert property (property_n78) else $error("property_n78 not held! ");
property_n79_assert : assert property (property_n79) else $error("property_n79 not held! ");
property_n80_assert : assert property (property_n80) else $error("property_n80 not held! ");
property_n81_assert : assert property (property_n81) else $error("property_n81 not held! ");
property_n82_assert : assert property (property_n82) else $error("property_n82 not held! ");
property_n83_assert : assert property (property_n83) else $error("property_n83 not held! ");
property_n84_assert : assert property (property_n84) else $error("property_n84 not held! ");
property_n85_assert : assert property (property_n85) else $error("property_n85 not held! ");
property_n86_assert : assert property (property_n86) else $error("property_n86 not held! ");
property_n87_assert : assert property (property_n87) else $error("property_n87 not held! ");
property_n88_assert : assert property (property_n88) else $error("property_n88 not held! ");
property_n89_assert : assert property (property_n89) else $error("property_n89 not held! ");
property_n90_assert : assert property (property_n90) else $error("property_n90 not held! ");
property_n91_assert : assert property (property_n91) else $error("property_n91 not held! ");
property_n92_assert : assert property (property_n92) else $error("property_n92 not held! ");
property_n93_assert : assert property (property_n93) else $error("property_n93 not held! ");
property_n94_assert : assert property (property_n94) else $error("property_n94 not held! ");
property_n95_assert : assert property (property_n95) else $error("property_n95 not held! ");
property_n96_assert : assert property (property_n96) else $error("property_n96 not held! ");
property_n97_assert : assert property (property_n97) else $error("property_n97 not held! ");
property_n98_assert : assert property (property_n98) else $error("property_n98 not held! ");
property_n99_assert : assert property (property_n99) else $error("property_n99 not held! ");
property_n100_assert : assert property (property_n100) else $error("property_n100 not held! ");
property_n101_assert : assert property (property_n101) else $error("property_n101 not held! ");
property_n102_assert : assert property (property_n102) else $error("property_n102 not held! ");
property_n103_assert : assert property (property_n103) else $error("property_n103 not held! ");
property_n104_assert : assert property (property_n104) else $error("property_n104 not held! ");
property_n105_assert : assert property (property_n105) else $error("property_n105 not held! ");
property_n106_assert : assert property (property_n106) else $error("property_n106 not held! ");
property_n107_assert : assert property (property_n107) else $error("property_n107 not held! ");
property_n108_assert : assert property (property_n108) else $error("property_n108 not held! ");
property_n109_assert : assert property (property_n109) else $error("property_n109 not held! ");
property_n110_assert : assert property (property_n110) else $error("property_n110 not held! ");
property_n111_assert : assert property (property_n111) else $error("property_n111 not held! ");
property_n112_assert : assert property (property_n112) else $error("property_n112 not held! ");
property_n113_assert : assert property (property_n113) else $error("property_n113 not held! ");
property_n114_assert : assert property (property_n114) else $error("property_n114 not held! ");
property_n115_assert : assert property (property_n115) else $error("property_n115 not held! ");
property_n116_assert : assert property (property_n116) else $error("property_n116 not held! ");
property_n117_assert : assert property (property_n117) else $error("property_n117 not held! ");
property_n118_assert : assert property (property_n118) else $error("property_n118 not held! ");
property_n119_assert : assert property (property_n119) else $error("property_n119 not held! ");
property_n120_assert : assert property (property_n120) else $error("property_n120 not held! ");
property_n121_assert : assert property (property_n121) else $error("property_n121 not held! ");
property_n122_assert : assert property (property_n122) else $error("property_n122 not held! ");
property_n123_assert : assert property (property_n123) else $error("property_n123 not held! ");
property_n124_assert : assert property (property_n124) else $error("property_n124 not held! ");
property_n125_assert : assert property (property_n125) else $error("property_n125 not held! ");
property_n126_assert : assert property (property_n126) else $error("property_n126 not held! ");
property_n127_assert : assert property (property_n127) else $error("property_n127 not held! ");
property_n128_assert : assert property (property_n128) else $error("property_n128 not held! ");
property_n129_assert : assert property (property_n129) else $error("property_n129 not held! ");
property_n130_assert : assert property (property_n130) else $error("property_n130 not held! ");
property_n131_assert : assert property (property_n131) else $error("property_n131 not held! ");
property_n132_assert : assert property (property_n132) else $error("property_n132 not held! ");
property_n133_assert : assert property (property_n133) else $error("property_n133 not held! ");
property_n134_assert : assert property (property_n134) else $error("property_n134 not held! ");
property_n135_assert : assert property (property_n135) else $error("property_n135 not held! ");
property_n136_assert : assert property (property_n136) else $error("property_n136 not held! ");
property_n137_assert : assert property (property_n137) else $error("property_n137 not held! ");
property_n138_assert : assert property (property_n138) else $error("property_n138 not held! ");
property_n139_assert : assert property (property_n139) else $error("property_n139 not held! ");
property_n140_assert : assert property (property_n140) else $error("property_n140 not held! ");
property_n141_assert : assert property (property_n141) else $error("property_n141 not held! ");
property_n142_assert : assert property (property_n142) else $error("property_n142 not held! ");
property_n143_assert : assert property (property_n143) else $error("property_n143 not held! ");
property_n144_assert : assert property (property_n144) else $error("property_n144 not held! ");
property_n145_assert : assert property (property_n145) else $error("property_n145 not held! ");
property_n146_assert : assert property (property_n146) else $error("property_n146 not held! ");
property_n147_assert : assert property (property_n147) else $error("property_n147 not held! ");
property_n148_assert : assert property (property_n148) else $error("property_n148 not held! ");
property_n149_assert : assert property (property_n149) else $error("property_n149 not held! ");
property_n150_assert : assert property (property_n150) else $error("property_n150 not held! ");
property_n151_assert : assert property (property_n151) else $error("property_n151 not held! ");
property_n152_assert : assert property (property_n152) else $error("property_n152 not held! ");
property_n153_assert : assert property (property_n153) else $error("property_n153 not held! ");
property_n154_assert : assert property (property_n154) else $error("property_n154 not held! ");
property_n155_assert : assert property (property_n155) else $error("property_n155 not held! ");
property_n156_assert : assert property (property_n156) else $error("property_n156 not held! ");
property_n157_assert : assert property (property_n157) else $error("property_n157 not held! ");
property_n158_assert : assert property (property_n158) else $error("property_n158 not held! ");
property_n159_assert : assert property (property_n159) else $error("property_n159 not held! ");
property_n160_assert : assert property (property_n160) else $error("property_n160 not held! ");
property_n161_assert : assert property (property_n161) else $error("property_n161 not held! ");
property_n162_assert : assert property (property_n162) else $error("property_n162 not held! ");
property_n163_assert : assert property (property_n163) else $error("property_n163 not held! ");
property_n164_assert : assert property (property_n164) else $error("property_n164 not held! ");
property_n165_assert : assert property (property_n165) else $error("property_n165 not held! ");
property_n166_assert : assert property (property_n166) else $error("property_n166 not held! ");
property_n167_assert : assert property (property_n167) else $error("property_n167 not held! ");
property_n168_assert : assert property (property_n168) else $error("property_n168 not held! ");
property_n169_assert : assert property (property_n169) else $error("property_n169 not held! ");
property_n170_assert : assert property (property_n170) else $error("property_n170 not held! ");
property_n171_assert : assert property (property_n171) else $error("property_n171 not held! ");
property_n172_assert : assert property (property_n172) else $error("property_n172 not held! ");
property_n173_assert : assert property (property_n173) else $error("property_n173 not held! ");
property_n174_assert : assert property (property_n174) else $error("property_n174 not held! ");
property_n175_assert : assert property (property_n175) else $error("property_n175 not held! ");
property_n176_assert : assert property (property_n176) else $error("property_n176 not held! ");
property_n177_assert : assert property (property_n177) else $error("property_n177 not held! ");
property_n178_assert : assert property (property_n178) else $error("property_n178 not held! ");
property_n179_assert : assert property (property_n179) else $error("property_n179 not held! ");
property_n180_assert : assert property (property_n180) else $error("property_n180 not held! ");
property_n181_assert : assert property (property_n181) else $error("property_n181 not held! ");
property_n182_assert : assert property (property_n182) else $error("property_n182 not held! ");
property_n183_assert : assert property (property_n183) else $error("property_n183 not held! ");
property_n184_assert : assert property (property_n184) else $error("property_n184 not held! ");
property_n185_assert : assert property (property_n185) else $error("property_n185 not held! ");
property_n186_assert : assert property (property_n186) else $error("property_n186 not held! ");
property_n187_assert : assert property (property_n187) else $error("property_n187 not held! ");
property_n188_assert : assert property (property_n188) else $error("property_n188 not held! ");
property_n189_assert : assert property (property_n189) else $error("property_n189 not held! ");
property_n190_assert : assert property (property_n190) else $error("property_n190 not held! ");
property_n191_assert : assert property (property_n191) else $error("property_n191 not held! ");
property_n192_assert : assert property (property_n192) else $error("property_n192 not held! ");
property_n193_assert : assert property (property_n193) else $error("property_n193 not held! ");
property_n194_assert : assert property (property_n194) else $error("property_n194 not held! ");
property_n195_assert : assert property (property_n195) else $error("property_n195 not held! ");
property_n196_assert : assert property (property_n196) else $error("property_n196 not held! ");
property_n197_assert : assert property (property_n197) else $error("property_n197 not held! ");
property_n198_assert : assert property (property_n198) else $error("property_n198 not held! ");
property_n199_assert : assert property (property_n199) else $error("property_n199 not held! ");
property_n200_assert : assert property (property_n200) else $error("property_n200 not held! ");
property_n201_assert : assert property (property_n201) else $error("property_n201 not held! ");
property_n202_assert : assert property (property_n202) else $error("property_n202 not held! ");
property_n203_assert : assert property (property_n203) else $error("property_n203 not held! ");
property_n204_assert : assert property (property_n204) else $error("property_n204 not held! ");
property_n205_assert : assert property (property_n205) else $error("property_n205 not held! ");
property_n206_assert : assert property (property_n206) else $error("property_n206 not held! ");
property_n207_assert : assert property (property_n207) else $error("property_n207 not held! ");
property_n208_assert : assert property (property_n208) else $error("property_n208 not held! ");
property_n209_assert : assert property (property_n209) else $error("property_n209 not held! ");
property_n210_assert : assert property (property_n210) else $error("property_n210 not held! ");
property_n211_assert : assert property (property_n211) else $error("property_n211 not held! ");
property_n212_assert : assert property (property_n212) else $error("property_n212 not held! ");
property_n213_assert : assert property (property_n213) else $error("property_n213 not held! ");
property_n214_assert : assert property (property_n214) else $error("property_n214 not held! ");
property_n215_assert : assert property (property_n215) else $error("property_n215 not held! ");
property_n216_assert : assert property (property_n216) else $error("property_n216 not held! ");
property_n217_assert : assert property (property_n217) else $error("property_n217 not held! ");
property_n218_assert : assert property (property_n218) else $error("property_n218 not held! ");
property_n219_assert : assert property (property_n219) else $error("property_n219 not held! ");
property_n220_assert : assert property (property_n220) else $error("property_n220 not held! ");
property_n221_assert : assert property (property_n221) else $error("property_n221 not held! ");
property_n222_assert : assert property (property_n222) else $error("property_n222 not held! ");
property_n223_assert : assert property (property_n223) else $error("property_n223 not held! ");
property_n224_assert : assert property (property_n224) else $error("property_n224 not held! ");
property_n225_assert : assert property (property_n225) else $error("property_n225 not held! ");
property_n226_assert : assert property (property_n226) else $error("property_n226 not held! ");
property_n227_assert : assert property (property_n227) else $error("property_n227 not held! ");
property_n228_assert : assert property (property_n228) else $error("property_n228 not held! ");
property_n229_assert : assert property (property_n229) else $error("property_n229 not held! ");
property_n230_assert : assert property (property_n230) else $error("property_n230 not held! ");
property_n231_assert : assert property (property_n231) else $error("property_n231 not held! ");
property_n232_assert : assert property (property_n232) else $error("property_n232 not held! ");
property_n233_assert : assert property (property_n233) else $error("property_n233 not held! ");
property_n234_assert : assert property (property_n234) else $error("property_n234 not held! ");
property_n235_assert : assert property (property_n235) else $error("property_n235 not held! ");
property_n236_assert : assert property (property_n236) else $error("property_n236 not held! ");
property_n237_assert : assert property (property_n237) else $error("property_n237 not held! ");
property_n238_assert : assert property (property_n238) else $error("property_n238 not held! ");
property_n239_assert : assert property (property_n239) else $error("property_n239 not held! ");
property_n240_assert : assert property (property_n240) else $error("property_n240 not held! ");
property_n241_assert : assert property (property_n241) else $error("property_n241 not held! ");
property_n242_assert : assert property (property_n242) else $error("property_n242 not held! ");
property_n243_assert : assert property (property_n243) else $error("property_n243 not held! ");
property_n244_assert : assert property (property_n244) else $error("property_n244 not held! ");
property_n248_assert : assert property (property_n248) else $error("property_n248 not held! ");
property_n249_assert : assert property (property_n249) else $error("property_n249 not held! ");
property_n251_assert : assert property (property_n251) else $error("property_n251 not held! ");
property_n252_assert : assert property (property_n252) else $error("property_n252 not held! ");
property_n256_assert : assert property (property_n256) else $error("property_n256 not held! ");
property_n258_assert : assert property (property_n258) else $error("property_n258 not held! ");
property_n260_assert : assert property (property_n260) else $error("property_n260 not held! ");
property_n261_assert : assert property (property_n261) else $error("property_n261 not held! ");
property_n264_assert : assert property (property_n264) else $error("property_n264 not held! ");
property_n265_assert : assert property (property_n265) else $error("property_n265 not held! ");

property_n279_assert : assert property (property_n279) else $error("property_n279 not held! ");

property_n281_assert : assert property (property_n281) else $error("property_n281 not held! ");

property_n285_assert : assert property (property_n285) else $error("property_n285 not held! ");

property_n287_assert : assert property (property_n287) else $error("property_n287 not held! ");

property_n289_assert : assert property (property_n289) else $error("property_n289 not held! ");
property_n290_assert : assert property (property_n290) else $error("property_n290 not held! ");
property_n291_assert : assert property (property_n291) else $error("property_n291 not held! ");
property_n292_assert : assert property (property_n292) else $error("property_n292 not held! ");
property_n293_assert : assert property (property_n293) else $error("property_n293 not held! ");
property_n294_assert : assert property (property_n294) else $error("property_n294 not held! ");
property_n295_assert : assert property (property_n295) else $error("property_n295 not held! ");
property_n296_assert : assert property (property_n296) else $error("property_n296 not held! ");
property_n297_assert : assert property (property_n297) else $error("property_n297 not held! ");
property_n298_assert : assert property (property_n298) else $error("property_n298 not held! ");
property_n299_assert : assert property (property_n299) else $error("property_n299 not held! ");
property_n300_assert : assert property (property_n300) else $error("property_n300 not held! ");

property_n305_assert : assert property (property_n305) else $error("property_n305 not held! ");

property_n311_assert : assert property (property_n311) else $error("property_n311 not held! ");
property_n312_assert : assert property (property_n312) else $error("property_n312 not held! ");
property_n313_assert : assert property (property_n313) else $error("property_n313 not held! ");
property_n316_assert : assert property (property_n316) else $error("property_n316 not held! ");
property_n317_assert : assert property (property_n317) else $error("property_n317 not held! ");
property_n318_assert : assert property (property_n318) else $error("property_n318 not held! ");
property_n322_assert : assert property (property_n322) else $error("property_n322 not held! ");
property_n323_assert : assert property (property_n323) else $error("property_n323 not held! ");
property_n324_assert : assert property (property_n324) else $error("property_n324 not held! ");
property_n325_assert : assert property (property_n325) else $error("property_n325 not held! ");
property_n327_assert : assert property (property_n327) else $error("property_n327 not held! ");
property_n328_assert : assert property (property_n328) else $error("property_n328 not held! ");
property_n342_assert : assert property (property_n342) else $error("property_n342 not held! ");
property_n344_assert : assert property (property_n344) else $error("property_n344 not held! ");
property_n345_assert : assert property (property_n345) else $error("property_n345 not held! ");
property_n347_assert : assert property (property_n347) else $error("property_n347 not held! ");
property_n348_assert : assert property (property_n348) else $error("property_n348 not held! ");
property_n354_assert : assert property (property_n354) else $error("property_n354 not held! ");
property_n357_assert : assert property (property_n357) else $error("property_n357 not held! ");
property_n358_assert : assert property (property_n358) else $error("property_n358 not held! ");
property_n359_assert : assert property (property_n359) else $error("property_n359 not held! ");
property_n360_assert : assert property (property_n360) else $error("property_n360 not held! ");
property_n361_assert : assert property (property_n361) else $error("property_n361 not held! ");
property_n362_assert : assert property (property_n362) else $error("property_n362 not held! ");
property_n363_assert : assert property (property_n363) else $error("property_n363 not held! ");
property_n366_assert : assert property (property_n366) else $error("property_n366 not held! ");
property_n367_assert : assert property (property_n367) else $error("property_n367 not held! ");
property_n369_assert : assert property (property_n369) else $error("property_n369 not held! ");
property_n370_assert : assert property (property_n370) else $error("property_n370 not held! ");
property_n371_assert : assert property (property_n371) else $error("property_n371 not held! ");
property_n372_assert : assert property (property_n372) else $error("property_n372 not held! ");
property_n373_assert : assert property (property_n373) else $error("property_n373 not held! ");
property_n374_assert : assert property (property_n374) else $error("property_n374 not held! ");
property_n377_assert : assert property (property_n377) else $error("property_n377 not held! ");
property_n378_assert : assert property (property_n378) else $error("property_n378 not held! ");
property_n379_assert : assert property (property_n379) else $error("property_n379 not held! ");
property_n381_assert : assert property (property_n381) else $error("property_n381 not held! ");
property_n382_assert : assert property (property_n382) else $error("property_n382 not held! ");
property_n383_assert : assert property (property_n383) else $error("property_n383 not held! ");
property_n385_assert : assert property (property_n385) else $error("property_n385 not held! ");
property_n387_assert : assert property (property_n387) else $error("property_n387 not held! ");
property_n388_assert : assert property (property_n388) else $error("property_n388 not held! ");
property_n391_assert : assert property (property_n391) else $error("property_n391 not held! ");
property_n393_assert : assert property (property_n393) else $error("property_n393 not held! ");
property_n394_assert : assert property (property_n394) else $error("property_n394 not held! ");
property_n395_assert : assert property (property_n395) else $error("property_n395 not held! ");
property_n396_assert : assert property (property_n396) else $error("property_n396 not held! ");
property_n398_assert : assert property (property_n398) else $error("property_n398 not held! ");
property_n399_assert : assert property (property_n399) else $error("property_n399 not held! ");
property_n401_assert : assert property (property_n401) else $error("property_n401 not held! ");
property_n402_assert : assert property (property_n402) else $error("property_n402 not held! ");
property_n403_assert : assert property (property_n403) else $error("property_n403 not held! ");
property_n404_assert : assert property (property_n404) else $error("property_n404 not held! ");
property_n405_assert : assert property (property_n405) else $error("property_n405 not held! ");
property_n406_assert : assert property (property_n406) else $error("property_n406 not held! ");
property_n407_assert : assert property (property_n407) else $error("property_n407 not held! ");
property_n408_assert : assert property (property_n408) else $error("property_n408 not held! ");
property_n409_assert : assert property (property_n409) else $error("property_n409 not held! ");
property_n410_assert : assert property (property_n410) else $error("property_n410 not held! ");
property_n411_assert : assert property (property_n411) else $error("property_n411 not held! ");
property_n412_assert : assert property (property_n412) else $error("property_n412 not held! ");
property_n413_assert : assert property (property_n413) else $error("property_n413 not held! ");
property_n414_assert : assert property (property_n414) else $error("property_n414 not held! ");
property_n415_assert : assert property (property_n415) else $error("property_n415 not held! ");
property_n416_assert : assert property (property_n416) else $error("property_n416 not held! ");
property_n417_assert : assert property (property_n417) else $error("property_n417 not held! ");
property_n418_assert : assert property (property_n418) else $error("property_n418 not held! ");
property_n419_assert : assert property (property_n419) else $error("property_n419 not held! ");
property_n420_assert : assert property (property_n420) else $error("property_n420 not held! ");
property_n421_assert : assert property (property_n421) else $error("property_n421 not held! ");
property_n422_assert : assert property (property_n422) else $error("property_n422 not held! ");
property_n423_assert : assert property (property_n423) else $error("property_n423 not held! ");
property_n424_assert : assert property (property_n424) else $error("property_n424 not held! ");
property_n425_assert : assert property (property_n425) else $error("property_n425 not held! ");
property_n428_assert : assert property (property_n428) else $error("property_n428 not held! ");
property_n431_assert : assert property (property_n431) else $error("property_n431 not held! ");
property_n432_assert : assert property (property_n432) else $error("property_n432 not held! ");
property_n435_assert : assert property (property_n435) else $error("property_n435 not held! ");
property_n436_assert : assert property (property_n436) else $error("property_n436 not held! ");
property_n437_assert : assert property (property_n437) else $error("property_n437 not held! ");
property_n438_assert : assert property (property_n438) else $error("property_n438 not held! ");
property_n439_assert : assert property (property_n439) else $error("property_n439 not held! ");
property_n440_assert : assert property (property_n440) else $error("property_n440 not held! ");
property_n441_assert : assert property (property_n441) else $error("property_n441 not held! ");
property_n442_assert : assert property (property_n442) else $error("property_n442 not held! ");
property_n443_assert : assert property (property_n443) else $error("property_n443 not held! ");
property_n444_assert : assert property (property_n444) else $error("property_n444 not held! ");
property_n445_assert : assert property (property_n445) else $error("property_n445 not held! ");
property_n446_assert : assert property (property_n446) else $error("property_n446 not held! ");
property_n447_assert : assert property (property_n447) else $error("property_n447 not held! ");
property_n448_assert : assert property (property_n448) else $error("property_n448 not held! ");
property_n449_assert : assert property (property_n449) else $error("property_n449 not held! ");
property_n450_assert : assert property (property_n450) else $error("property_n450 not held! ");
property_n451_assert : assert property (property_n451) else $error("property_n451 not held! ");
property_n453_assert : assert property (property_n453) else $error("property_n453 not held! ");
property_n454_assert : assert property (property_n454) else $error("property_n454 not held! ");
property_n455_assert : assert property (property_n455) else $error("property_n455 not held! ");
property_n456_assert : assert property (property_n456) else $error("property_n456 not held! ");
property_n457_assert : assert property (property_n457) else $error("property_n457 not held! ");
property_n458_assert : assert property (property_n458) else $error("property_n458 not held! ");
property_n459_assert : assert property (property_n459) else $error("property_n459 not held! ");
property_n460_assert : assert property (property_n460) else $error("property_n460 not held! ");
property_n461_assert : assert property (property_n461) else $error("property_n461 not held! ");
property_n462_assert : assert property (property_n462) else $error("property_n462 not held! ");
property_n463_assert : assert property (property_n463) else $error("property_n463 not held! ");
property_n464_assert : assert property (property_n464) else $error("property_n464 not held! ");
property_n465_assert : assert property (property_n465) else $error("property_n465 not held! ");
property_n466_assert : assert property (property_n466) else $error("property_n466 not held! ");
property_n467_assert : assert property (property_n467) else $error("property_n467 not held! ");
property_n469_assert : assert property (property_n469) else $error("property_n469 not held! ");
property_n470_assert : assert property (property_n470) else $error("property_n470 not held! ");
property_n471_assert : assert property (property_n471) else $error("property_n471 not held! ");
property_n473_assert : assert property (property_n473) else $error("property_n473 not held! ");
property_n474_assert : assert property (property_n474) else $error("property_n474 not held! ");
property_n475_assert : assert property (property_n475) else $error("property_n475 not held! ");
property_n476_assert : assert property (property_n476) else $error("property_n476 not held! ");
property_n477_assert : assert property (property_n477) else $error("property_n477 not held! ");
property_n478_assert : assert property (property_n478) else $error("property_n478 not held! ");
property_n480_assert : assert property (property_n480) else $error("property_n480 not held! ");
property_n482_assert : assert property (property_n482) else $error("property_n482 not held! ");
property_n483_assert : assert property (property_n483) else $error("property_n483 not held! ");
property_n484_assert : assert property (property_n484) else $error("property_n484 not held! ");
property_n486_assert : assert property (property_n486) else $error("property_n486 not held! ");
property_n487_assert : assert property (property_n487) else $error("property_n487 not held! ");
property_n488_assert : assert property (property_n488) else $error("property_n488 not held! ");
property_n489_assert : assert property (property_n489) else $error("property_n489 not held! ");

  
endmodule
